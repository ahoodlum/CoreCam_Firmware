library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

---- Uncomment the following library declaration if instantiating
---- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity datarom is
    Port ( CLK : in std_logic;
           ADDR : in std_logic_vector(19 DOWNTO 0);
           DOUT : out std_logic_vector(35 DOWNTO 0)
           );
end datarom;


architecture behavior of datarom is

begin 

main : process (CLK)
begin    
if (falling_edge(CLK)) then 
    case ADDR is

		when x"00000" => DOUT <= x"0000001a1";
		when x"00001" => DOUT <= x"000000120";
		when x"00002" => DOUT <= x"000200141";
		when x"00003" => DOUT <= x"000200140";
		when x"00004" => DOUT <= x"000001121";
		when x"00005" => DOUT <= x"0000011a0";
		when x"00006" => DOUT <= x"0002011c1";
		when x"00007" => DOUT <= x"0002011c0";
		when x"00008" => DOUT <= x"0000001a1";
		when x"00009" => DOUT <= x"000000120";
		when x"0000a" => DOUT <= x"000200141";
		when x"0000b" => DOUT <= x"000200140";
		when x"0000c" => DOUT <= x"000001121";
		when x"0000d" => DOUT <= x"0000011a0";
		when x"0000e" => DOUT <= x"0002011c1";
		when x"0000f" => DOUT <= x"0002011c0";
		when x"00010" => DOUT <= x"0000021a1";
		when x"00011" => DOUT <= x"000002120";
		when x"00012" => DOUT <= x"000202141";
		when x"00013" => DOUT <= x"000202140";
		when x"00014" => DOUT <= x"000003121";
		when x"00015" => DOUT <= x"0000031a0";
		when x"00016" => DOUT <= x"0002031c1";
		when x"00017" => DOUT <= x"0002031c0";
		when x"00018" => DOUT <= x"0000021a1";
		when x"00019" => DOUT <= x"000002120";
		when x"0001a" => DOUT <= x"000202141";
		when x"0001b" => DOUT <= x"000202140";
		when x"0001c" => DOUT <= x"000003121";
		when x"0001d" => DOUT <= x"0000031a0";
		when x"0001e" => DOUT <= x"0002031c1";
		when x"0001f" => DOUT <= x"0002031c0";
		when x"00020" => DOUT <= x"0000021a1";
		when x"00021" => DOUT <= x"000002120";
		when x"00022" => DOUT <= x"000202141";
		when x"00023" => DOUT <= x"000202140";
		when x"00024" => DOUT <= x"000003121";
		when x"00025" => DOUT <= x"0000031a0";
		when x"00026" => DOUT <= x"0002031c1";
		when x"00027" => DOUT <= x"0002031c0";
		when x"00028" => DOUT <= x"0000021a1";
		when x"00029" => DOUT <= x"000002120";
		when x"0002a" => DOUT <= x"000202141";
		when x"0002b" => DOUT <= x"000202140";
		when x"0002c" => DOUT <= x"000003121";
		when x"0002d" => DOUT <= x"0000031a0";
		when x"0002e" => DOUT <= x"0002031c1";
		when x"0002f" => DOUT <= x"0002031c0";
		when x"00030" => DOUT <= x"0000021a1";
		when x"00031" => DOUT <= x"000002120";
		when x"00032" => DOUT <= x"000202141";
		when x"00033" => DOUT <= x"000202140";
		when x"00034" => DOUT <= x"000003121";
		when x"00035" => DOUT <= x"0000031a0";
		when x"00036" => DOUT <= x"0002031c1";
		when x"00037" => DOUT <= x"0002031c0";
		when x"00038" => DOUT <= x"0000021a1";
		when x"00039" => DOUT <= x"000002120";
		when x"0003a" => DOUT <= x"000202141";
		when x"0003b" => DOUT <= x"000202140";
		when x"0003c" => DOUT <= x"000003121";
		when x"0003d" => DOUT <= x"0000031a0";
		when x"0003e" => DOUT <= x"0002031c1";
		when x"0003f" => DOUT <= x"0002031c0";
		when x"00040" => DOUT <= x"0000021a1";
		when x"00041" => DOUT <= x"000002120";
		when x"00042" => DOUT <= x"000202141";
		when x"00043" => DOUT <= x"000202140";
		when x"00044" => DOUT <= x"000003121";
		when x"00045" => DOUT <= x"0000031a0";
		when x"00046" => DOUT <= x"0002031c1";
		when x"00047" => DOUT <= x"0002031c0";
		when x"00048" => DOUT <= x"0000021a1";
		when x"00049" => DOUT <= x"000002120";
		when x"0004a" => DOUT <= x"000202141";
		when x"0004b" => DOUT <= x"000202140";
		when x"0004c" => DOUT <= x"000003121";
		when x"0004d" => DOUT <= x"0000031a0";
		when x"0004e" => DOUT <= x"0002031c1";
		when x"0004f" => DOUT <= x"0002031c0";
		when x"00050" => DOUT <= x"0000021a1";
		when x"00051" => DOUT <= x"000002120";
		when x"00052" => DOUT <= x"000202141";
		when x"00053" => DOUT <= x"000202140";
		when x"00054" => DOUT <= x"000003121";
		when x"00055" => DOUT <= x"0000031a0";
		when x"00056" => DOUT <= x"0002031c1";
		when x"00057" => DOUT <= x"0002031c0";
		when x"00058" => DOUT <= x"0000021a1";
		when x"00059" => DOUT <= x"000002120";
		when x"0005a" => DOUT <= x"000202141";
		when x"0005b" => DOUT <= x"000202140";
		when x"0005c" => DOUT <= x"000003121";
		when x"0005d" => DOUT <= x"0000031a0";
		when x"0005e" => DOUT <= x"0002031c1";
		when x"0005f" => DOUT <= x"0002031c0";
		when x"00060" => DOUT <= x"0000021a1";
		when x"00061" => DOUT <= x"000002120";
		when x"00062" => DOUT <= x"000202141";
		when x"00063" => DOUT <= x"000202140";
		when x"00064" => DOUT <= x"000003121";
		when x"00065" => DOUT <= x"0000031a0";
		when x"00066" => DOUT <= x"0002031c1";
		when x"00067" => DOUT <= x"0002031c0";
		when x"00068" => DOUT <= x"0000021a1";
		when x"00069" => DOUT <= x"000002120";
		when x"0006a" => DOUT <= x"000202141";
		when x"0006b" => DOUT <= x"000202140";
		when x"0006c" => DOUT <= x"000003121";
		when x"0006d" => DOUT <= x"0000031a0";
		when x"0006e" => DOUT <= x"0002031c1";
		when x"0006f" => DOUT <= x"0002031c0";
		when x"00070" => DOUT <= x"0000021a1";
		when x"00071" => DOUT <= x"000002120";
		when x"00072" => DOUT <= x"000202141";
		when x"00073" => DOUT <= x"000202140";
		when x"00074" => DOUT <= x"000003121";
		when x"00075" => DOUT <= x"0000031a0";
		when x"00076" => DOUT <= x"0002031c1";
		when x"00077" => DOUT <= x"0002031c0";
		when x"00078" => DOUT <= x"0000021a1";
		when x"00079" => DOUT <= x"000002120";
		when x"0007a" => DOUT <= x"000202141";
		when x"0007b" => DOUT <= x"000202140";
		when x"0007c" => DOUT <= x"000003121";
		when x"0007d" => DOUT <= x"0000031a0";
		when x"0007e" => DOUT <= x"0002031c1";
		when x"0007f" => DOUT <= x"0002031c0";
		when x"00080" => DOUT <= x"0000021a1";
		when x"00081" => DOUT <= x"000002120";
		when x"00082" => DOUT <= x"000202141";
		when x"00083" => DOUT <= x"000202140";
		when x"00084" => DOUT <= x"000003121";
		when x"00085" => DOUT <= x"0000031a0";
		when x"00086" => DOUT <= x"0002031c1";
		when x"00087" => DOUT <= x"0002031c0";
		when x"00088" => DOUT <= x"0000021a1";
		when x"00089" => DOUT <= x"000002120";
		when x"0008a" => DOUT <= x"000202141";
		when x"0008b" => DOUT <= x"000202140";
		when x"0008c" => DOUT <= x"000003121";
		when x"0008d" => DOUT <= x"0000031a0";
		when x"0008e" => DOUT <= x"0002031c1";
		when x"0008f" => DOUT <= x"0002031c0";
		when x"00090" => DOUT <= x"0000021a1";
		when x"00091" => DOUT <= x"000002120";
		when x"00092" => DOUT <= x"000202141";
		when x"00093" => DOUT <= x"000202140";
		when x"00094" => DOUT <= x"000003121";
		when x"00095" => DOUT <= x"0000031a0";
		when x"00096" => DOUT <= x"0002031c1";
		when x"00097" => DOUT <= x"0002031c0";
		when x"00098" => DOUT <= x"0000021a1";
		when x"00099" => DOUT <= x"000002120";
		when x"0009a" => DOUT <= x"000202141";
		when x"0009b" => DOUT <= x"000202140";
		when x"0009c" => DOUT <= x"000003121";
		when x"0009d" => DOUT <= x"0000031a0";
		when x"0009e" => DOUT <= x"0002031c1";
		when x"0009f" => DOUT <= x"0002031c0";
		when x"000a0" => DOUT <= x"0000021a1";
		when x"000a1" => DOUT <= x"000002120";
		when x"000a2" => DOUT <= x"000202141";
		when x"000a3" => DOUT <= x"000202140";
		when x"000a4" => DOUT <= x"000003121";
		when x"000a5" => DOUT <= x"0000031a0";
		when x"000a6" => DOUT <= x"0002031c1";
		when x"000a7" => DOUT <= x"0002031c0";
		when x"000a8" => DOUT <= x"0000021a1";
		when x"000a9" => DOUT <= x"000002120";
		when x"000aa" => DOUT <= x"000202141";
		when x"000ab" => DOUT <= x"000202140";
		when x"000ac" => DOUT <= x"000003121";
		when x"000ad" => DOUT <= x"0000031a0";
		when x"000ae" => DOUT <= x"0002031c1";
		when x"000af" => DOUT <= x"0002031c0";
		when x"000b0" => DOUT <= x"0000021a1";
		when x"000b1" => DOUT <= x"000002120";
		when x"000b2" => DOUT <= x"000202141";
		when x"000b3" => DOUT <= x"000202140";
		when x"000b4" => DOUT <= x"000003121";
		when x"000b5" => DOUT <= x"0000031a0";
		when x"000b6" => DOUT <= x"0002031c1";
		when x"000b7" => DOUT <= x"0002031c0";
		when x"000b8" => DOUT <= x"0000021a1";
		when x"000b9" => DOUT <= x"000002120";
		when x"000ba" => DOUT <= x"000202141";
		when x"000bb" => DOUT <= x"000202140";
		when x"000bc" => DOUT <= x"000003121";
		when x"000bd" => DOUT <= x"0000031a0";
		when x"000be" => DOUT <= x"0002031c1";
		when x"000bf" => DOUT <= x"0002031c0";
		when x"000c0" => DOUT <= x"0000021a1";
		when x"000c1" => DOUT <= x"000002120";
		when x"000c2" => DOUT <= x"000202141";
		when x"000c3" => DOUT <= x"000202140";
		when x"000c4" => DOUT <= x"000003121";
		when x"000c5" => DOUT <= x"0000031a0";
		when x"000c6" => DOUT <= x"0002031c1";
		when x"000c7" => DOUT <= x"0002031c0";
		when x"000c8" => DOUT <= x"0000021a1";
		when x"000c9" => DOUT <= x"000002120";
		when x"000ca" => DOUT <= x"000202141";
		when x"000cb" => DOUT <= x"000202140";
		when x"000cc" => DOUT <= x"000003121";
		when x"000cd" => DOUT <= x"0000031a0";
		when x"000ce" => DOUT <= x"0002031c1";
		when x"000cf" => DOUT <= x"0002031c0";
		when x"000d0" => DOUT <= x"0000021a1";
		when x"000d1" => DOUT <= x"000002120";
		when x"000d2" => DOUT <= x"000202141";
		when x"000d3" => DOUT <= x"000202140";
		when x"000d4" => DOUT <= x"000003121";
		when x"000d5" => DOUT <= x"0000031a0";
		when x"000d6" => DOUT <= x"0002031c1";
		when x"000d7" => DOUT <= x"0002031c0";
		when x"000d8" => DOUT <= x"0000021a1";
		when x"000d9" => DOUT <= x"000002120";
		when x"000da" => DOUT <= x"000202141";
		when x"000db" => DOUT <= x"000202140";
		when x"000dc" => DOUT <= x"000003121";
		when x"000dd" => DOUT <= x"0000031a0";
		when x"000de" => DOUT <= x"0002031c1";
		when x"000df" => DOUT <= x"0002031c0";
		when x"000e0" => DOUT <= x"0000021a1";
		when x"000e1" => DOUT <= x"000002120";
		when x"000e2" => DOUT <= x"000202141";
		when x"000e3" => DOUT <= x"000202140";
		when x"000e4" => DOUT <= x"000003121";
		when x"000e5" => DOUT <= x"0000031a0";
		when x"000e6" => DOUT <= x"0002031c1";
		when x"000e7" => DOUT <= x"0002031c0";
		when x"000e8" => DOUT <= x"0000021a1";
		when x"000e9" => DOUT <= x"000002120";
		when x"000ea" => DOUT <= x"000202141";
		when x"000eb" => DOUT <= x"000202140";
		when x"000ec" => DOUT <= x"000003121";
		when x"000ed" => DOUT <= x"0000031a0";
		when x"000ee" => DOUT <= x"0002031c1";
		when x"000ef" => DOUT <= x"0002031c0";
		when x"000f0" => DOUT <= x"0000021a1";
		when x"000f1" => DOUT <= x"000002120";
		when x"000f2" => DOUT <= x"000202141";
		when x"000f3" => DOUT <= x"000202140";
		when x"000f4" => DOUT <= x"000003121";
		when x"000f5" => DOUT <= x"0000031a0";
		when x"000f6" => DOUT <= x"0002031c1";
		when x"000f7" => DOUT <= x"0002031c0";
		when x"000f8" => DOUT <= x"0000021a1";
		when x"000f9" => DOUT <= x"000002120";
		when x"000fa" => DOUT <= x"000202141";
		when x"000fb" => DOUT <= x"000202140";
		when x"000fc" => DOUT <= x"000003121";
		when x"000fd" => DOUT <= x"0000031a0";
		when x"000fe" => DOUT <= x"0002031c1";
		when x"000ff" => DOUT <= x"0002031c0";
		when x"00100" => DOUT <= x"0000021a1";
		when x"00101" => DOUT <= x"000002120";
		when x"00102" => DOUT <= x"000202141";
		when x"00103" => DOUT <= x"000202140";
		when x"00104" => DOUT <= x"000003121";
		when x"00105" => DOUT <= x"0000031a0";
		when x"00106" => DOUT <= x"0002031c1";
		when x"00107" => DOUT <= x"0002031c0";
		when x"00108" => DOUT <= x"0000021a1";
		when x"00109" => DOUT <= x"000002120";
		when x"0010a" => DOUT <= x"000202141";
		when x"0010b" => DOUT <= x"000202140";
		when x"0010c" => DOUT <= x"000003121";
		when x"0010d" => DOUT <= x"0000031a0";
		when x"0010e" => DOUT <= x"0002031c1";
		when x"0010f" => DOUT <= x"0002031c0";
		when x"00110" => DOUT <= x"0000021a1";
		when x"00111" => DOUT <= x"000002120";
		when x"00112" => DOUT <= x"000202141";
		when x"00113" => DOUT <= x"000202140";
		when x"00114" => DOUT <= x"000003121";
		when x"00115" => DOUT <= x"0000031a0";
		when x"00116" => DOUT <= x"0002031c1";
		when x"00117" => DOUT <= x"0002031c0";
		when x"00118" => DOUT <= x"0000021a1";
		when x"00119" => DOUT <= x"000002120";
		when x"0011a" => DOUT <= x"000202141";
		when x"0011b" => DOUT <= x"000202140";
		when x"0011c" => DOUT <= x"000003121";
		when x"0011d" => DOUT <= x"0000031a0";
		when x"0011e" => DOUT <= x"0002031c1";
		when x"0011f" => DOUT <= x"0002031c0";
		when x"00120" => DOUT <= x"0000021a1";
		when x"00121" => DOUT <= x"000002120";
		when x"00122" => DOUT <= x"000202141";
		when x"00123" => DOUT <= x"000202140";
		when x"00124" => DOUT <= x"000003121";
		when x"00125" => DOUT <= x"0000031a0";
		when x"00126" => DOUT <= x"0002031c1";
		when x"00127" => DOUT <= x"0002031c0";
		when x"00128" => DOUT <= x"0000021a1";
		when x"00129" => DOUT <= x"000002120";
		when x"0012a" => DOUT <= x"000202141";
		when x"0012b" => DOUT <= x"000202140";
		when x"0012c" => DOUT <= x"000003121";
		when x"0012d" => DOUT <= x"0000031a0";
		when x"0012e" => DOUT <= x"0002031c1";
		when x"0012f" => DOUT <= x"0002031c0";
		when x"00130" => DOUT <= x"0000021a1";
		when x"00131" => DOUT <= x"000002120";
		when x"00132" => DOUT <= x"000202141";
		when x"00133" => DOUT <= x"000202140";
		when x"00134" => DOUT <= x"000003121";
		when x"00135" => DOUT <= x"0000031a0";
		when x"00136" => DOUT <= x"0002031c1";
		when x"00137" => DOUT <= x"0002031c0";
		when x"00138" => DOUT <= x"0000021a1";
		when x"00139" => DOUT <= x"000002120";
		when x"0013a" => DOUT <= x"000202141";
		when x"0013b" => DOUT <= x"000202140";
		when x"0013c" => DOUT <= x"000003121";
		when x"0013d" => DOUT <= x"0000031a0";
		when x"0013e" => DOUT <= x"0002031c1";
		when x"0013f" => DOUT <= x"0002031c0";
		when x"00140" => DOUT <= x"0000021a1";
		when x"00141" => DOUT <= x"000002120";
		when x"00142" => DOUT <= x"000202141";
		when x"00143" => DOUT <= x"000202140";
		when x"00144" => DOUT <= x"000003121";
		when x"00145" => DOUT <= x"0000031a0";
		when x"00146" => DOUT <= x"0002031c1";
		when x"00147" => DOUT <= x"0002031c0";
		when x"00148" => DOUT <= x"0000021a1";
		when x"00149" => DOUT <= x"000002120";
		when x"0014a" => DOUT <= x"000202141";
		when x"0014b" => DOUT <= x"000202140";
		when x"0014c" => DOUT <= x"000003121";
		when x"0014d" => DOUT <= x"0000031a0";
		when x"0014e" => DOUT <= x"0002031c1";
		when x"0014f" => DOUT <= x"0002031c0";
		when x"00150" => DOUT <= x"0000021a1";
		when x"00151" => DOUT <= x"000002120";
		when x"00152" => DOUT <= x"000202141";
		when x"00153" => DOUT <= x"000202140";
		when x"00154" => DOUT <= x"000003121";
		when x"00155" => DOUT <= x"0000031a0";
		when x"00156" => DOUT <= x"0002031c1";
		when x"00157" => DOUT <= x"0002031c0";
		when x"00158" => DOUT <= x"0000021a1";
		when x"00159" => DOUT <= x"000002120";
		when x"0015a" => DOUT <= x"000202141";
		when x"0015b" => DOUT <= x"000202140";
		when x"0015c" => DOUT <= x"000003121";
		when x"0015d" => DOUT <= x"0000031a0";
		when x"0015e" => DOUT <= x"0002031c1";
		when x"0015f" => DOUT <= x"0002031c0";
		when x"00160" => DOUT <= x"0000021a1";
		when x"00161" => DOUT <= x"000002120";
		when x"00162" => DOUT <= x"000202141";
		when x"00163" => DOUT <= x"000202140";
		when x"00164" => DOUT <= x"000003121";
		when x"00165" => DOUT <= x"0000031a0";
		when x"00166" => DOUT <= x"0002031c1";
		when x"00167" => DOUT <= x"0002031c0";
		when x"00168" => DOUT <= x"0000021a1";
		when x"00169" => DOUT <= x"000002120";
		when x"0016a" => DOUT <= x"000202141";
		when x"0016b" => DOUT <= x"000202140";
		when x"0016c" => DOUT <= x"000003121";
		when x"0016d" => DOUT <= x"0000031a0";
		when x"0016e" => DOUT <= x"0002031c1";
		when x"0016f" => DOUT <= x"0002031c0";
		when x"00170" => DOUT <= x"0000021a1";
		when x"00171" => DOUT <= x"000002120";
		when x"00172" => DOUT <= x"000202141";
		when x"00173" => DOUT <= x"000202140";
		when x"00174" => DOUT <= x"000003121";
		when x"00175" => DOUT <= x"0000031a0";
		when x"00176" => DOUT <= x"0002031c1";
		when x"00177" => DOUT <= x"0002031c0";
		when x"00178" => DOUT <= x"0000021a1";
		when x"00179" => DOUT <= x"000002120";
		when x"0017a" => DOUT <= x"000202141";
		when x"0017b" => DOUT <= x"000202140";
		when x"0017c" => DOUT <= x"000003121";
		when x"0017d" => DOUT <= x"0000031a0";
		when x"0017e" => DOUT <= x"0002031c1";
		when x"0017f" => DOUT <= x"0002031c0";
		when x"00180" => DOUT <= x"0000021a1";
		when x"00181" => DOUT <= x"000002120";
		when x"00182" => DOUT <= x"000202141";
		when x"00183" => DOUT <= x"000202140";
		when x"00184" => DOUT <= x"000003121";
		when x"00185" => DOUT <= x"0000031a0";
		when x"00186" => DOUT <= x"0002031c1";
		when x"00187" => DOUT <= x"0002031c0";
		when x"00188" => DOUT <= x"0000021a1";
		when x"00189" => DOUT <= x"000002120";
		when x"0018a" => DOUT <= x"000202141";
		when x"0018b" => DOUT <= x"000202140";
		when x"0018c" => DOUT <= x"000003121";
		when x"0018d" => DOUT <= x"0000031a0";
		when x"0018e" => DOUT <= x"0002031c1";
		when x"0018f" => DOUT <= x"0002031c0";
		when x"00190" => DOUT <= x"0000021a1";
		when x"00191" => DOUT <= x"000002120";
		when x"00192" => DOUT <= x"000202141";
		when x"00193" => DOUT <= x"000202140";
		when x"00194" => DOUT <= x"000003121";
		when x"00195" => DOUT <= x"0000031a0";
		when x"00196" => DOUT <= x"0002031c1";
		when x"00197" => DOUT <= x"0002031c0";
		when x"00198" => DOUT <= x"0000021a1";
		when x"00199" => DOUT <= x"000002120";
		when x"0019a" => DOUT <= x"000202141";
		when x"0019b" => DOUT <= x"000202140";
		when x"0019c" => DOUT <= x"000003121";
		when x"0019d" => DOUT <= x"0000031a0";
		when x"0019e" => DOUT <= x"0002031c1";
		when x"0019f" => DOUT <= x"0002031c0";
		when x"001a0" => DOUT <= x"0000021a1";
		when x"001a1" => DOUT <= x"000002120";
		when x"001a2" => DOUT <= x"000202141";
		when x"001a3" => DOUT <= x"000202140";
		when x"001a4" => DOUT <= x"000003121";
		when x"001a5" => DOUT <= x"0000031a0";
		when x"001a6" => DOUT <= x"0002031c1";
		when x"001a7" => DOUT <= x"0002031c0";
		when x"001a8" => DOUT <= x"0000021a1";
		when x"001a9" => DOUT <= x"000002120";
		when x"001aa" => DOUT <= x"000202141";
		when x"001ab" => DOUT <= x"000202140";
		when x"001ac" => DOUT <= x"000003121";
		when x"001ad" => DOUT <= x"0000031a0";
		when x"001ae" => DOUT <= x"0002031c1";
		when x"001af" => DOUT <= x"0002031c0";
		when x"001b0" => DOUT <= x"0000021a1";
		when x"001b1" => DOUT <= x"000002120";
		when x"001b2" => DOUT <= x"000202141";
		when x"001b3" => DOUT <= x"000202140";
		when x"001b4" => DOUT <= x"000003121";
		when x"001b5" => DOUT <= x"0000031a0";
		when x"001b6" => DOUT <= x"0002031c1";
		when x"001b7" => DOUT <= x"0002031c0";
		when x"001b8" => DOUT <= x"0000021a1";
		when x"001b9" => DOUT <= x"000002120";
		when x"001ba" => DOUT <= x"000202141";
		when x"001bb" => DOUT <= x"000202140";
		when x"001bc" => DOUT <= x"000003121";
		when x"001bd" => DOUT <= x"0000031a0";
		when x"001be" => DOUT <= x"0002031c1";
		when x"001bf" => DOUT <= x"0002031c0";
		when x"001c0" => DOUT <= x"0000021a1";
		when x"001c1" => DOUT <= x"000002120";
		when x"001c2" => DOUT <= x"000202141";
		when x"001c3" => DOUT <= x"000202140";
		when x"001c4" => DOUT <= x"000003121";
		when x"001c5" => DOUT <= x"0000031a0";
		when x"001c6" => DOUT <= x"0002031c1";
		when x"001c7" => DOUT <= x"0002031c0";
		when x"001c8" => DOUT <= x"0000021a1";
		when x"001c9" => DOUT <= x"000002120";
		when x"001ca" => DOUT <= x"000202141";
		when x"001cb" => DOUT <= x"000202140";
		when x"001cc" => DOUT <= x"000003121";
		when x"001cd" => DOUT <= x"0000031a0";
		when x"001ce" => DOUT <= x"0002031c1";
		when x"001cf" => DOUT <= x"0002031c0";
		when x"001d0" => DOUT <= x"0000021a1";
		when x"001d1" => DOUT <= x"000002120";
		when x"001d2" => DOUT <= x"000202141";
		when x"001d3" => DOUT <= x"000202140";
		when x"001d4" => DOUT <= x"000003121";
		when x"001d5" => DOUT <= x"0000031a0";
		when x"001d6" => DOUT <= x"0002031c1";
		when x"001d7" => DOUT <= x"0002031c0";
		when x"001d8" => DOUT <= x"0000021a1";
		when x"001d9" => DOUT <= x"000002120";
		when x"001da" => DOUT <= x"000202141";
		when x"001db" => DOUT <= x"000202140";
		when x"001dc" => DOUT <= x"000003121";
		when x"001dd" => DOUT <= x"0000031a0";
		when x"001de" => DOUT <= x"0002031c1";
		when x"001df" => DOUT <= x"0002031c0";
		when x"001e0" => DOUT <= x"0000021a1";
		when x"001e1" => DOUT <= x"000002120";
		when x"001e2" => DOUT <= x"000202141";
		when x"001e3" => DOUT <= x"000202140";
		when x"001e4" => DOUT <= x"000003121";
		when x"001e5" => DOUT <= x"0000031a0";
		when x"001e6" => DOUT <= x"0002031c1";
		when x"001e7" => DOUT <= x"0002031c0";
		when x"001e8" => DOUT <= x"0000021a1";
		when x"001e9" => DOUT <= x"000002120";
		when x"001ea" => DOUT <= x"000202141";
		when x"001eb" => DOUT <= x"000202140";
		when x"001ec" => DOUT <= x"000003121";
		when x"001ed" => DOUT <= x"0000031a0";
		when x"001ee" => DOUT <= x"0002031c1";
		when x"001ef" => DOUT <= x"0002031c0";
		when x"001f0" => DOUT <= x"0000021a1";
		when x"001f1" => DOUT <= x"000002120";
		when x"001f2" => DOUT <= x"000202141";
		when x"001f3" => DOUT <= x"000202140";
		when x"001f4" => DOUT <= x"000003121";
		when x"001f5" => DOUT <= x"0000031a0";
		when x"001f6" => DOUT <= x"0002031c1";
		when x"001f7" => DOUT <= x"0002031c0";
		when x"001f8" => DOUT <= x"0000021a1";
		when x"001f9" => DOUT <= x"000002120";
		when x"001fa" => DOUT <= x"000202141";
		when x"001fb" => DOUT <= x"000202140";
		when x"001fc" => DOUT <= x"000003121";
		when x"001fd" => DOUT <= x"0000031a0";
		when x"001fe" => DOUT <= x"0002031c1";
		when x"001ff" => DOUT <= x"0002031c0";
		when x"00200" => DOUT <= x"0000021a1";
		when x"00201" => DOUT <= x"000002120";
		when x"00202" => DOUT <= x"000202141";
		when x"00203" => DOUT <= x"000202140";
		when x"00204" => DOUT <= x"000003121";
		when x"00205" => DOUT <= x"0000031a0";
		when x"00206" => DOUT <= x"0002031c1";
		when x"00207" => DOUT <= x"0002031c0";
		when x"00208" => DOUT <= x"0000021a1";
		when x"00209" => DOUT <= x"000002120";
		when x"0020a" => DOUT <= x"000202141";
		when x"0020b" => DOUT <= x"000202140";
		when x"0020c" => DOUT <= x"000003121";
		when x"0020d" => DOUT <= x"0000031a0";
		when x"0020e" => DOUT <= x"0002031c1";
		when x"0020f" => DOUT <= x"0002031c0";
		when x"00210" => DOUT <= x"0000021a1";
		when x"00211" => DOUT <= x"000002120";
		when x"00212" => DOUT <= x"000202141";
		when x"00213" => DOUT <= x"000202140";
		when x"00214" => DOUT <= x"000003121";
		when x"00215" => DOUT <= x"0000031a0";
		when x"00216" => DOUT <= x"0002031c1";
		when x"00217" => DOUT <= x"0002031c0";
		when x"00218" => DOUT <= x"0000021a1";
		when x"00219" => DOUT <= x"000002120";
		when x"0021a" => DOUT <= x"000202141";
		when x"0021b" => DOUT <= x"000202140";
		when x"0021c" => DOUT <= x"000003121";
		when x"0021d" => DOUT <= x"0000031a0";
		when x"0021e" => DOUT <= x"0002031c1";
		when x"0021f" => DOUT <= x"0002031c0";
		when x"00220" => DOUT <= x"0000021a1";
		when x"00221" => DOUT <= x"000002120";
		when x"00222" => DOUT <= x"000202141";
		when x"00223" => DOUT <= x"000202140";
		when x"00224" => DOUT <= x"000003121";
		when x"00225" => DOUT <= x"0000031a0";
		when x"00226" => DOUT <= x"0002031c1";
		when x"00227" => DOUT <= x"0002031c0";
		when x"00228" => DOUT <= x"0000021a1";
		when x"00229" => DOUT <= x"000002120";
		when x"0022a" => DOUT <= x"000202141";
		when x"0022b" => DOUT <= x"000202140";
		when x"0022c" => DOUT <= x"000003121";
		when x"0022d" => DOUT <= x"0000031a0";
		when x"0022e" => DOUT <= x"0002031c1";
		when x"0022f" => DOUT <= x"0002031c0";
		when x"00230" => DOUT <= x"0000021a1";
		when x"00231" => DOUT <= x"000002120";
		when x"00232" => DOUT <= x"000202141";
		when x"00233" => DOUT <= x"000202140";
		when x"00234" => DOUT <= x"000003121";
		when x"00235" => DOUT <= x"0000031a0";
		when x"00236" => DOUT <= x"0002031c1";
		when x"00237" => DOUT <= x"0002031c0";
		when x"00238" => DOUT <= x"0000021a1";
		when x"00239" => DOUT <= x"000002120";
		when x"0023a" => DOUT <= x"000202141";
		when x"0023b" => DOUT <= x"000202140";
		when x"0023c" => DOUT <= x"000003121";
		when x"0023d" => DOUT <= x"0000031a0";
		when x"0023e" => DOUT <= x"0002031c1";
		when x"0023f" => DOUT <= x"0002031c0";
		when x"00240" => DOUT <= x"0000021a1";
		when x"00241" => DOUT <= x"000002120";
		when x"00242" => DOUT <= x"000202141";
		when x"00243" => DOUT <= x"000202140";
		when x"00244" => DOUT <= x"000003121";
		when x"00245" => DOUT <= x"0000031a0";
		when x"00246" => DOUT <= x"0002031c1";
		when x"00247" => DOUT <= x"0002031c0";
		when x"00248" => DOUT <= x"0000021a1";
		when x"00249" => DOUT <= x"000002120";
		when x"0024a" => DOUT <= x"000202141";
		when x"0024b" => DOUT <= x"000202140";
		when x"0024c" => DOUT <= x"000003121";
		when x"0024d" => DOUT <= x"0000031a0";
		when x"0024e" => DOUT <= x"0002031c1";
		when x"0024f" => DOUT <= x"0002031c0";
		when x"00250" => DOUT <= x"0000021a1";
		when x"00251" => DOUT <= x"000002120";
		when x"00252" => DOUT <= x"000202141";
		when x"00253" => DOUT <= x"000202140";
		when x"00254" => DOUT <= x"000003121";
		when x"00255" => DOUT <= x"0000031a0";
		when x"00256" => DOUT <= x"0002031c1";
		when x"00257" => DOUT <= x"0002031c0";
		when x"00258" => DOUT <= x"0000021a1";
		when x"00259" => DOUT <= x"000002120";
		when x"0025a" => DOUT <= x"000202141";
		when x"0025b" => DOUT <= x"000202140";
		when x"0025c" => DOUT <= x"000003121";
		when x"0025d" => DOUT <= x"0000031a0";
		when x"0025e" => DOUT <= x"0002031c1";
		when x"0025f" => DOUT <= x"0002031c0";
		when x"00260" => DOUT <= x"0000021a1";
		when x"00261" => DOUT <= x"000002120";
		when x"00262" => DOUT <= x"000202141";
		when x"00263" => DOUT <= x"000202140";
		when x"00264" => DOUT <= x"000003121";
		when x"00265" => DOUT <= x"0000031a0";
		when x"00266" => DOUT <= x"0002031c1";
		when x"00267" => DOUT <= x"0002031c0";
		when x"00268" => DOUT <= x"0000021a1";
		when x"00269" => DOUT <= x"000002120";
		when x"0026a" => DOUT <= x"000202141";
		when x"0026b" => DOUT <= x"000202140";
		when x"0026c" => DOUT <= x"000003121";
		when x"0026d" => DOUT <= x"0000031a0";
		when x"0026e" => DOUT <= x"0002031c1";
		when x"0026f" => DOUT <= x"0002031c0";
		when x"00270" => DOUT <= x"0000021a1";
		when x"00271" => DOUT <= x"000002120";
		when x"00272" => DOUT <= x"000202141";
		when x"00273" => DOUT <= x"000202140";
		when x"00274" => DOUT <= x"000003121";
		when x"00275" => DOUT <= x"0000031a0";
		when x"00276" => DOUT <= x"0002031c1";
		when x"00277" => DOUT <= x"0002031c0";
		when x"00278" => DOUT <= x"0000021a1";
		when x"00279" => DOUT <= x"000002120";
		when x"0027a" => DOUT <= x"000202141";
		when x"0027b" => DOUT <= x"000202140";
		when x"0027c" => DOUT <= x"000003121";
		when x"0027d" => DOUT <= x"0000031a0";
		when x"0027e" => DOUT <= x"0002031c1";
		when x"0027f" => DOUT <= x"0002031c0";
		when x"00280" => DOUT <= x"0000021a1";
		when x"00281" => DOUT <= x"000002120";
		when x"00282" => DOUT <= x"000202141";
		when x"00283" => DOUT <= x"000202140";
		when x"00284" => DOUT <= x"000003121";
		when x"00285" => DOUT <= x"0000031a0";
		when x"00286" => DOUT <= x"0002031c1";
		when x"00287" => DOUT <= x"0002031c0";
		when x"00288" => DOUT <= x"0000021a1";
		when x"00289" => DOUT <= x"000002120";
		when x"0028a" => DOUT <= x"000202141";
		when x"0028b" => DOUT <= x"000202140";
		when x"0028c" => DOUT <= x"000003121";
		when x"0028d" => DOUT <= x"0000031a0";
		when x"0028e" => DOUT <= x"0002031c1";
		when x"0028f" => DOUT <= x"0002031c0";
		when x"00290" => DOUT <= x"0000021a1";
		when x"00291" => DOUT <= x"000002120";
		when x"00292" => DOUT <= x"000202141";
		when x"00293" => DOUT <= x"000202140";
		when x"00294" => DOUT <= x"000003121";
		when x"00295" => DOUT <= x"0000031a0";
		when x"00296" => DOUT <= x"0002031c1";
		when x"00297" => DOUT <= x"0002031c0";
		when x"00298" => DOUT <= x"0000021a1";
		when x"00299" => DOUT <= x"000002120";
		when x"0029a" => DOUT <= x"000202141";
		when x"0029b" => DOUT <= x"000202140";
		when x"0029c" => DOUT <= x"000003121";
		when x"0029d" => DOUT <= x"0000031a0";
		when x"0029e" => DOUT <= x"0002031c1";
		when x"0029f" => DOUT <= x"0002031c0";
		when x"002a0" => DOUT <= x"0000021a1";
		when x"002a1" => DOUT <= x"000002120";
		when x"002a2" => DOUT <= x"000202141";
		when x"002a3" => DOUT <= x"000202140";
		when x"002a4" => DOUT <= x"000003121";
		when x"002a5" => DOUT <= x"0000031a0";
		when x"002a6" => DOUT <= x"0002031c1";
		when x"002a7" => DOUT <= x"0002031c0";
		when x"002a8" => DOUT <= x"0000021a1";
		when x"002a9" => DOUT <= x"000002120";
		when x"002aa" => DOUT <= x"000202141";
		when x"002ab" => DOUT <= x"000202140";
		when x"002ac" => DOUT <= x"000003121";
		when x"002ad" => DOUT <= x"0000031a0";
		when x"002ae" => DOUT <= x"0002031c1";
		when x"002af" => DOUT <= x"0002031c0";
		when x"002b0" => DOUT <= x"0000021a1";
		when x"002b1" => DOUT <= x"000002120";
		when x"002b2" => DOUT <= x"000202141";
		when x"002b3" => DOUT <= x"000202140";
		when x"002b4" => DOUT <= x"000003121";
		when x"002b5" => DOUT <= x"0000031a0";
		when x"002b6" => DOUT <= x"0002031c1";
		when x"002b7" => DOUT <= x"0002031c0";
		when x"002b8" => DOUT <= x"0000021a1";
		when x"002b9" => DOUT <= x"000002120";
		when x"002ba" => DOUT <= x"000202141";
		when x"002bb" => DOUT <= x"000202140";
		when x"002bc" => DOUT <= x"000003121";
		when x"002bd" => DOUT <= x"0000031a0";
		when x"002be" => DOUT <= x"0002031c1";
		when x"002bf" => DOUT <= x"0002031c0";
		when x"002c0" => DOUT <= x"0000021a1";
		when x"002c1" => DOUT <= x"000002120";
		when x"002c2" => DOUT <= x"000202141";
		when x"002c3" => DOUT <= x"000202140";
		when x"002c4" => DOUT <= x"000003121";
		when x"002c5" => DOUT <= x"0000031a0";
		when x"002c6" => DOUT <= x"0002031c1";
		when x"002c7" => DOUT <= x"0002031c0";
		when x"002c8" => DOUT <= x"0000021a1";
		when x"002c9" => DOUT <= x"000002120";
		when x"002ca" => DOUT <= x"000202141";
		when x"002cb" => DOUT <= x"000202140";
		when x"002cc" => DOUT <= x"000003121";
		when x"002cd" => DOUT <= x"0000031a0";
		when x"002ce" => DOUT <= x"0002031c1";
		when x"002cf" => DOUT <= x"0002031c0";
		when x"002d0" => DOUT <= x"0000021a1";
		when x"002d1" => DOUT <= x"000002120";
		when x"002d2" => DOUT <= x"000202141";
		when x"002d3" => DOUT <= x"000202140";
		when x"002d4" => DOUT <= x"000003121";
		when x"002d5" => DOUT <= x"0000031a0";
		when x"002d6" => DOUT <= x"0002031c1";
		when x"002d7" => DOUT <= x"0002031c0";
		when x"002d8" => DOUT <= x"0000021a1";
		when x"002d9" => DOUT <= x"000002120";
		when x"002da" => DOUT <= x"000202141";
		when x"002db" => DOUT <= x"000202140";
		when x"002dc" => DOUT <= x"000003121";
		when x"002dd" => DOUT <= x"0000031a0";
		when x"002de" => DOUT <= x"0002031c1";
		when x"002df" => DOUT <= x"0002031c0";
		when x"002e0" => DOUT <= x"0000021a1";
		when x"002e1" => DOUT <= x"000002120";
		when x"002e2" => DOUT <= x"000202141";
		when x"002e3" => DOUT <= x"000202140";
		when x"002e4" => DOUT <= x"000003121";
		when x"002e5" => DOUT <= x"0000031a0";
		when x"002e6" => DOUT <= x"0002031c1";
		when x"002e7" => DOUT <= x"0002031c0";
		when x"002e8" => DOUT <= x"0000021a1";
		when x"002e9" => DOUT <= x"000002120";
		when x"002ea" => DOUT <= x"000202141";
		when x"002eb" => DOUT <= x"000202140";
		when x"002ec" => DOUT <= x"000003121";
		when x"002ed" => DOUT <= x"0000031a0";
		when x"002ee" => DOUT <= x"0002031c1";
		when x"002ef" => DOUT <= x"0002031c0";
		when x"002f0" => DOUT <= x"0000021a1";
		when x"002f1" => DOUT <= x"000002120";
		when x"002f2" => DOUT <= x"000202141";
		when x"002f3" => DOUT <= x"000202140";
		when x"002f4" => DOUT <= x"000003121";
		when x"002f5" => DOUT <= x"0000031a0";
		when x"002f6" => DOUT <= x"0002031c1";
		when x"002f7" => DOUT <= x"0002031c0";
		when x"002f8" => DOUT <= x"0000021a1";
		when x"002f9" => DOUT <= x"000002120";
		when x"002fa" => DOUT <= x"000202141";
		when x"002fb" => DOUT <= x"000202140";
		when x"002fc" => DOUT <= x"000003121";
		when x"002fd" => DOUT <= x"0000031a0";
		when x"002fe" => DOUT <= x"0002031c1";
		when x"002ff" => DOUT <= x"0002031c0";
		when x"00300" => DOUT <= x"0000021a1";
		when x"00301" => DOUT <= x"000002120";
		when x"00302" => DOUT <= x"000202141";
		when x"00303" => DOUT <= x"000202140";
		when x"00304" => DOUT <= x"000003121";
		when x"00305" => DOUT <= x"0000031a0";
		when x"00306" => DOUT <= x"0002031c1";
		when x"00307" => DOUT <= x"0002031c0";
		when x"00308" => DOUT <= x"0000021a1";
		when x"00309" => DOUT <= x"000002120";
		when x"0030a" => DOUT <= x"000202141";
		when x"0030b" => DOUT <= x"000202140";
		when x"0030c" => DOUT <= x"000003121";
		when x"0030d" => DOUT <= x"0000031a0";
		when x"0030e" => DOUT <= x"0002031c1";
		when x"0030f" => DOUT <= x"0002031c0";
		when x"00310" => DOUT <= x"0000021a1";
		when x"00311" => DOUT <= x"000002120";
		when x"00312" => DOUT <= x"000202141";
		when x"00313" => DOUT <= x"000202140";
		when x"00314" => DOUT <= x"000003121";
		when x"00315" => DOUT <= x"0000031a0";
		when x"00316" => DOUT <= x"0002031c1";
		when x"00317" => DOUT <= x"0002031c0";
		when x"00318" => DOUT <= x"0000021a1";
		when x"00319" => DOUT <= x"000002120";
		when x"0031a" => DOUT <= x"000202141";
		when x"0031b" => DOUT <= x"000202140";
		when x"0031c" => DOUT <= x"000003121";
		when x"0031d" => DOUT <= x"0000031a0";
		when x"0031e" => DOUT <= x"0002031c1";
		when x"0031f" => DOUT <= x"0002031c0";
		when x"00320" => DOUT <= x"0000021a1";
		when x"00321" => DOUT <= x"000002120";
		when x"00322" => DOUT <= x"000202141";
		when x"00323" => DOUT <= x"000202140";
		when x"00324" => DOUT <= x"000003121";
		when x"00325" => DOUT <= x"0000031a0";
		when x"00326" => DOUT <= x"0002031c1";
		when x"00327" => DOUT <= x"0002031c0";
		when x"00328" => DOUT <= x"0000021a1";
		when x"00329" => DOUT <= x"000002120";
		when x"0032a" => DOUT <= x"000202141";
		when x"0032b" => DOUT <= x"000202140";
		when x"0032c" => DOUT <= x"000003121";
		when x"0032d" => DOUT <= x"0000031a0";
		when x"0032e" => DOUT <= x"0002031c1";
		when x"0032f" => DOUT <= x"0002031c0";
		when x"00330" => DOUT <= x"0000021a1";
		when x"00331" => DOUT <= x"000002120";
		when x"00332" => DOUT <= x"000202141";
		when x"00333" => DOUT <= x"000202140";
		when x"00334" => DOUT <= x"000003121";
		when x"00335" => DOUT <= x"0000031a0";
		when x"00336" => DOUT <= x"0002031c1";
		when x"00337" => DOUT <= x"0002031c0";
		when x"00338" => DOUT <= x"0000021a1";
		when x"00339" => DOUT <= x"000002120";
		when x"0033a" => DOUT <= x"000202141";
		when x"0033b" => DOUT <= x"000202140";
		when x"0033c" => DOUT <= x"000003121";
		when x"0033d" => DOUT <= x"0000031a0";
		when x"0033e" => DOUT <= x"0002031c1";
		when x"0033f" => DOUT <= x"0002031c0";
		when x"00340" => DOUT <= x"0000021a1";
		when x"00341" => DOUT <= x"000002120";
		when x"00342" => DOUT <= x"000202141";
		when x"00343" => DOUT <= x"000202140";
		when x"00344" => DOUT <= x"000003121";
		when x"00345" => DOUT <= x"0000031a0";
		when x"00346" => DOUT <= x"0002031c1";
		when x"00347" => DOUT <= x"0002031c0";
		when x"00348" => DOUT <= x"0000021a1";
		when x"00349" => DOUT <= x"000002120";
		when x"0034a" => DOUT <= x"000202141";
		when x"0034b" => DOUT <= x"000202140";
		when x"0034c" => DOUT <= x"000003121";
		when x"0034d" => DOUT <= x"0000031a0";
		when x"0034e" => DOUT <= x"0002031c1";
		when x"0034f" => DOUT <= x"0002031c0";
		when x"00350" => DOUT <= x"0000021a1";
		when x"00351" => DOUT <= x"000002120";
		when x"00352" => DOUT <= x"000202141";
		when x"00353" => DOUT <= x"000202140";
		when x"00354" => DOUT <= x"000003121";
		when x"00355" => DOUT <= x"0000031a0";
		when x"00356" => DOUT <= x"0002031c1";
		when x"00357" => DOUT <= x"0002031c0";
		when x"00358" => DOUT <= x"0000021a1";
		when x"00359" => DOUT <= x"000002120";
		when x"0035a" => DOUT <= x"000202141";
		when x"0035b" => DOUT <= x"000202140";
		when x"0035c" => DOUT <= x"000003121";
		when x"0035d" => DOUT <= x"0000031a0";
		when x"0035e" => DOUT <= x"0002031c1";
		when x"0035f" => DOUT <= x"0002031c0";
		when x"00360" => DOUT <= x"0000021a1";
		when x"00361" => DOUT <= x"000002120";
		when x"00362" => DOUT <= x"000202141";
		when x"00363" => DOUT <= x"000202140";
		when x"00364" => DOUT <= x"000003121";
		when x"00365" => DOUT <= x"0000031a0";
		when x"00366" => DOUT <= x"0002031c1";
		when x"00367" => DOUT <= x"0002031c0";
		when x"00368" => DOUT <= x"0000021a1";
		when x"00369" => DOUT <= x"000002120";
		when x"0036a" => DOUT <= x"000202141";
		when x"0036b" => DOUT <= x"000202140";
		when x"0036c" => DOUT <= x"000003121";
		when x"0036d" => DOUT <= x"0000031a0";
		when x"0036e" => DOUT <= x"0002031c1";
		when x"0036f" => DOUT <= x"0002031c0";
		when x"00370" => DOUT <= x"0000021a1";
		when x"00371" => DOUT <= x"000002120";
		when x"00372" => DOUT <= x"000202141";
		when x"00373" => DOUT <= x"000202140";
		when x"00374" => DOUT <= x"000003121";
		when x"00375" => DOUT <= x"0000031a0";
		when x"00376" => DOUT <= x"0002031c1";
		when x"00377" => DOUT <= x"0002031c0";
		when x"00378" => DOUT <= x"0000021a1";
		when x"00379" => DOUT <= x"000002120";
		when x"0037a" => DOUT <= x"000202141";
		when x"0037b" => DOUT <= x"000202140";
		when x"0037c" => DOUT <= x"000003121";
		when x"0037d" => DOUT <= x"0000031a0";
		when x"0037e" => DOUT <= x"0002031c1";
		when x"0037f" => DOUT <= x"0002031c0";
		when x"00380" => DOUT <= x"0000021a1";
		when x"00381" => DOUT <= x"000002120";
		when x"00382" => DOUT <= x"000202141";
		when x"00383" => DOUT <= x"000202140";
		when x"00384" => DOUT <= x"000003121";
		when x"00385" => DOUT <= x"0000031a0";
		when x"00386" => DOUT <= x"0002031c1";
		when x"00387" => DOUT <= x"0002031c0";
		when x"00388" => DOUT <= x"0000021a1";
		when x"00389" => DOUT <= x"000002120";
		when x"0038a" => DOUT <= x"000202141";
		when x"0038b" => DOUT <= x"000202140";
		when x"0038c" => DOUT <= x"000003121";
		when x"0038d" => DOUT <= x"0000031a0";
		when x"0038e" => DOUT <= x"0002031c1";
		when x"0038f" => DOUT <= x"0002031c0";
		when x"00390" => DOUT <= x"0000021a1";
		when x"00391" => DOUT <= x"000002120";
		when x"00392" => DOUT <= x"000202141";
		when x"00393" => DOUT <= x"000202140";
		when x"00394" => DOUT <= x"000003121";
		when x"00395" => DOUT <= x"0000031a0";
		when x"00396" => DOUT <= x"0002031c1";
		when x"00397" => DOUT <= x"0002031c0";
		when x"00398" => DOUT <= x"0000021a1";
		when x"00399" => DOUT <= x"000002120";
		when x"0039a" => DOUT <= x"000202141";
		when x"0039b" => DOUT <= x"000202140";
		when x"0039c" => DOUT <= x"000003121";
		when x"0039d" => DOUT <= x"0000031a0";
		when x"0039e" => DOUT <= x"0002031c1";
		when x"0039f" => DOUT <= x"0002031c0";
		when x"003a0" => DOUT <= x"0000021a1";
		when x"003a1" => DOUT <= x"000002120";
		when x"003a2" => DOUT <= x"000202141";
		when x"003a3" => DOUT <= x"000202140";
		when x"003a4" => DOUT <= x"000003121";
		when x"003a5" => DOUT <= x"0000031a0";
		when x"003a6" => DOUT <= x"0002031c1";
		when x"003a7" => DOUT <= x"0002031c0";
		when x"003a8" => DOUT <= x"0000021a1";
		when x"003a9" => DOUT <= x"000002120";
		when x"003aa" => DOUT <= x"000202141";
		when x"003ab" => DOUT <= x"000202140";
		when x"003ac" => DOUT <= x"000003121";
		when x"003ad" => DOUT <= x"0000031a0";
		when x"003ae" => DOUT <= x"0002031c1";
		when x"003af" => DOUT <= x"0002031c0";
		when x"003b0" => DOUT <= x"0000021a1";
		when x"003b1" => DOUT <= x"000002120";
		when x"003b2" => DOUT <= x"000202141";
		when x"003b3" => DOUT <= x"000202140";
		when x"003b4" => DOUT <= x"000003121";
		when x"003b5" => DOUT <= x"0000031a0";
		when x"003b6" => DOUT <= x"0002031c1";
		when x"003b7" => DOUT <= x"0002031c0";
		when x"003b8" => DOUT <= x"0000021a1";
		when x"003b9" => DOUT <= x"000002120";
		when x"003ba" => DOUT <= x"000202141";
		when x"003bb" => DOUT <= x"000202140";
		when x"003bc" => DOUT <= x"000003121";
		when x"003bd" => DOUT <= x"0000031a0";
		when x"003be" => DOUT <= x"0002031c1";
		when x"003bf" => DOUT <= x"0002031c0";
		when x"003c0" => DOUT <= x"0000021a1";
		when x"003c1" => DOUT <= x"000002120";
		when x"003c2" => DOUT <= x"000202141";
		when x"003c3" => DOUT <= x"000202140";
		when x"003c4" => DOUT <= x"000003121";
		when x"003c5" => DOUT <= x"0000031a0";
		when x"003c6" => DOUT <= x"0002031c1";
		when x"003c7" => DOUT <= x"0002031c0";
		when x"003c8" => DOUT <= x"0000021a1";
		when x"003c9" => DOUT <= x"000002120";
		when x"003ca" => DOUT <= x"000202141";
		when x"003cb" => DOUT <= x"000202140";
		when x"003cc" => DOUT <= x"000003121";
		when x"003cd" => DOUT <= x"0000031a0";
		when x"003ce" => DOUT <= x"0002031c1";
		when x"003cf" => DOUT <= x"0002031c0";
		when x"003d0" => DOUT <= x"0000021a1";
		when x"003d1" => DOUT <= x"000002120";
		when x"003d2" => DOUT <= x"000202141";
		when x"003d3" => DOUT <= x"000202140";
		when x"003d4" => DOUT <= x"000003121";
		when x"003d5" => DOUT <= x"0000031a0";
		when x"003d6" => DOUT <= x"0002031c1";
		when x"003d7" => DOUT <= x"0002031c0";
		when x"003d8" => DOUT <= x"0000021a1";
		when x"003d9" => DOUT <= x"000002120";
		when x"003da" => DOUT <= x"000202141";
		when x"003db" => DOUT <= x"000202140";
		when x"003dc" => DOUT <= x"000003121";
		when x"003dd" => DOUT <= x"0000031a0";
		when x"003de" => DOUT <= x"0002031c1";
		when x"003df" => DOUT <= x"0002031c0";
		when x"003e0" => DOUT <= x"0000021a1";
		when x"003e1" => DOUT <= x"000002120";
		when x"003e2" => DOUT <= x"000202141";
		when x"003e3" => DOUT <= x"000202140";
		when x"003e4" => DOUT <= x"000003121";
		when x"003e5" => DOUT <= x"0000031a0";
		when x"003e6" => DOUT <= x"0002031c1";
		when x"003e7" => DOUT <= x"0002031c0";
		when x"003e8" => DOUT <= x"0000021a1";
		when x"003e9" => DOUT <= x"000002120";
		when x"003ea" => DOUT <= x"000202141";
		when x"003eb" => DOUT <= x"000202140";
		when x"003ec" => DOUT <= x"000003121";
		when x"003ed" => DOUT <= x"0000031a0";
		when x"003ee" => DOUT <= x"0002031c1";
		when x"003ef" => DOUT <= x"0002031c0";
		when x"003f0" => DOUT <= x"0000021a1";
		when x"003f1" => DOUT <= x"000002120";
		when x"003f2" => DOUT <= x"000202141";
		when x"003f3" => DOUT <= x"000202140";
		when x"003f4" => DOUT <= x"000003121";
		when x"003f5" => DOUT <= x"0000031a0";
		when x"003f6" => DOUT <= x"0002031c1";
		when x"003f7" => DOUT <= x"0002031c0";
		when x"003f8" => DOUT <= x"0000021a1";
		when x"003f9" => DOUT <= x"000002120";
		when x"003fa" => DOUT <= x"000202141";
		when x"003fb" => DOUT <= x"000202140";
		when x"003fc" => DOUT <= x"000003121";
		when x"003fd" => DOUT <= x"0000031a0";
		when x"003fe" => DOUT <= x"0002031c1";
		when x"003ff" => DOUT <= x"0002031c0";
		when x"00400" => DOUT <= x"0000021a1";
		when x"00401" => DOUT <= x"000002120";
		when x"00402" => DOUT <= x"000202141";
		when x"00403" => DOUT <= x"000202140";
		when x"00404" => DOUT <= x"000003121";
		when x"00405" => DOUT <= x"0000031a0";
		when x"00406" => DOUT <= x"0002031c1";
		when x"00407" => DOUT <= x"0002031c0";
		when x"00408" => DOUT <= x"0000021a1";
		when x"00409" => DOUT <= x"000002120";
		when x"0040a" => DOUT <= x"000202141";
		when x"0040b" => DOUT <= x"000202140";
		when x"0040c" => DOUT <= x"000003121";
		when x"0040d" => DOUT <= x"0000031a0";
		when x"0040e" => DOUT <= x"0002031c1";
		when x"0040f" => DOUT <= x"0002031c0";
		when x"00410" => DOUT <= x"0000021a1";
		when x"00411" => DOUT <= x"000002120";
		when x"00412" => DOUT <= x"000202141";
		when x"00413" => DOUT <= x"000202140";
		when x"00414" => DOUT <= x"000003121";
		when x"00415" => DOUT <= x"0000031a0";
		when x"00416" => DOUT <= x"0002031c1";
		when x"00417" => DOUT <= x"0002031c0";
		when x"00418" => DOUT <= x"0000021a1";
		when x"00419" => DOUT <= x"000002120";
		when x"0041a" => DOUT <= x"000202141";
		when x"0041b" => DOUT <= x"000202140";
		when x"0041c" => DOUT <= x"000003121";
		when x"0041d" => DOUT <= x"0000031a0";
		when x"0041e" => DOUT <= x"0002031c1";
		when x"0041f" => DOUT <= x"0002031c0";
		when x"00420" => DOUT <= x"0000021a1";
		when x"00421" => DOUT <= x"000002120";
		when x"00422" => DOUT <= x"000202141";
		when x"00423" => DOUT <= x"000202140";
		when x"00424" => DOUT <= x"000003121";
		when x"00425" => DOUT <= x"0000031a0";
		when x"00426" => DOUT <= x"0002031c1";
		when x"00427" => DOUT <= x"0002031c0";
		when x"00428" => DOUT <= x"0000021a1";
		when x"00429" => DOUT <= x"000002120";
		when x"0042a" => DOUT <= x"000202141";
		when x"0042b" => DOUT <= x"000202140";
		when x"0042c" => DOUT <= x"000003121";
		when x"0042d" => DOUT <= x"0000031a0";
		when x"0042e" => DOUT <= x"0002031c1";
		when x"0042f" => DOUT <= x"0002031c0";
		when x"00430" => DOUT <= x"0000021a1";
		when x"00431" => DOUT <= x"000002120";
		when x"00432" => DOUT <= x"000202141";
		when x"00433" => DOUT <= x"000202140";
		when x"00434" => DOUT <= x"000003121";
		when x"00435" => DOUT <= x"0000031a0";
		when x"00436" => DOUT <= x"0002031c1";
		when x"00437" => DOUT <= x"0002031c0";
		when x"00438" => DOUT <= x"0000021a1";
		when x"00439" => DOUT <= x"000002120";
		when x"0043a" => DOUT <= x"000202141";
		when x"0043b" => DOUT <= x"000202140";
		when x"0043c" => DOUT <= x"000003121";
		when x"0043d" => DOUT <= x"0000031a0";
		when x"0043e" => DOUT <= x"0002031c1";
		when x"0043f" => DOUT <= x"0002031c0";
		when x"00440" => DOUT <= x"0000021a1";
		when x"00441" => DOUT <= x"000002120";
		when x"00442" => DOUT <= x"000202141";
		when x"00443" => DOUT <= x"000202140";
		when x"00444" => DOUT <= x"000003121";
		when x"00445" => DOUT <= x"0000031a0";
		when x"00446" => DOUT <= x"0002031c1";
		when x"00447" => DOUT <= x"0002031c0";
		when x"00448" => DOUT <= x"0000021a1";
		when x"00449" => DOUT <= x"000002120";
		when x"0044a" => DOUT <= x"000202141";
		when x"0044b" => DOUT <= x"000202140";
		when x"0044c" => DOUT <= x"000003121";
		when x"0044d" => DOUT <= x"0000031a0";
		when x"0044e" => DOUT <= x"0002031c1";
		when x"0044f" => DOUT <= x"0002031c0";
		when x"00450" => DOUT <= x"0000021a1";
		when x"00451" => DOUT <= x"000002120";
		when x"00452" => DOUT <= x"000202141";
		when x"00453" => DOUT <= x"000202140";
		when x"00454" => DOUT <= x"000003121";
		when x"00455" => DOUT <= x"0000031a0";
		when x"00456" => DOUT <= x"0002031c1";
		when x"00457" => DOUT <= x"0002031c0";
		when x"00458" => DOUT <= x"0000021a1";
		when x"00459" => DOUT <= x"000002120";
		when x"0045a" => DOUT <= x"000202141";
		when x"0045b" => DOUT <= x"000202140";
		when x"0045c" => DOUT <= x"000003121";
		when x"0045d" => DOUT <= x"0000031a0";
		when x"0045e" => DOUT <= x"0002031c1";
		when x"0045f" => DOUT <= x"0002031c0";
		when x"00460" => DOUT <= x"0000021a1";
		when x"00461" => DOUT <= x"000002120";
		when x"00462" => DOUT <= x"000202141";
		when x"00463" => DOUT <= x"000202140";
		when x"00464" => DOUT <= x"000003121";
		when x"00465" => DOUT <= x"0000031a0";
		when x"00466" => DOUT <= x"0002031c1";
		when x"00467" => DOUT <= x"0002031c0";
		when x"00468" => DOUT <= x"0000021a1";
		when x"00469" => DOUT <= x"000002120";
		when x"0046a" => DOUT <= x"000202141";
		when x"0046b" => DOUT <= x"000202140";
		when x"0046c" => DOUT <= x"000003121";
		when x"0046d" => DOUT <= x"0000031a0";
		when x"0046e" => DOUT <= x"0002031c1";
		when x"0046f" => DOUT <= x"0002031c0";
		when x"00470" => DOUT <= x"0000021a1";
		when x"00471" => DOUT <= x"000002120";
		when x"00472" => DOUT <= x"000202141";
		when x"00473" => DOUT <= x"000202140";
		when x"00474" => DOUT <= x"000003121";
		when x"00475" => DOUT <= x"0000031a0";
		when x"00476" => DOUT <= x"0002031c1";
		when x"00477" => DOUT <= x"0002031c0";
		when x"00478" => DOUT <= x"0000021a1";
		when x"00479" => DOUT <= x"000002120";
		when x"0047a" => DOUT <= x"000202141";
		when x"0047b" => DOUT <= x"000202140";
		when x"0047c" => DOUT <= x"000003121";
		when x"0047d" => DOUT <= x"0000031a0";
		when x"0047e" => DOUT <= x"0002031c1";
		when x"0047f" => DOUT <= x"0002031c0";
		when x"00480" => DOUT <= x"0000021a1";
		when x"00481" => DOUT <= x"000002120";
		when x"00482" => DOUT <= x"000202141";
		when x"00483" => DOUT <= x"000202140";
		when x"00484" => DOUT <= x"000003121";
		when x"00485" => DOUT <= x"0000031a0";
		when x"00486" => DOUT <= x"0002031c1";
		when x"00487" => DOUT <= x"0002031c0";
		when x"00488" => DOUT <= x"0000021a1";
		when x"00489" => DOUT <= x"000002120";
		when x"0048a" => DOUT <= x"000202141";
		when x"0048b" => DOUT <= x"000202140";
		when x"0048c" => DOUT <= x"000003121";
		when x"0048d" => DOUT <= x"0000031a0";
		when x"0048e" => DOUT <= x"0002031c1";
		when x"0048f" => DOUT <= x"0002031c0";
		when x"00490" => DOUT <= x"0000021a1";
		when x"00491" => DOUT <= x"000002120";
		when x"00492" => DOUT <= x"000202141";
		when x"00493" => DOUT <= x"000202140";
		when x"00494" => DOUT <= x"000003121";
		when x"00495" => DOUT <= x"0000031a0";
		when x"00496" => DOUT <= x"0002031c1";
		when x"00497" => DOUT <= x"0002031c0";
		when x"00498" => DOUT <= x"0000021a1";
		when x"00499" => DOUT <= x"000002120";
		when x"0049a" => DOUT <= x"000202141";
		when x"0049b" => DOUT <= x"000202140";
		when x"0049c" => DOUT <= x"000003121";
		when x"0049d" => DOUT <= x"0000031a0";
		when x"0049e" => DOUT <= x"0002031c1";
		when x"0049f" => DOUT <= x"0002031c0";
		when x"004a0" => DOUT <= x"0000021a1";
		when x"004a1" => DOUT <= x"000002120";
		when x"004a2" => DOUT <= x"000202141";
		when x"004a3" => DOUT <= x"000202140";
		when x"004a4" => DOUT <= x"000003121";
		when x"004a5" => DOUT <= x"0000031a0";
		when x"004a6" => DOUT <= x"0002031c1";
		when x"004a7" => DOUT <= x"0002031c0";
		when x"004a8" => DOUT <= x"0000021a1";
		when x"004a9" => DOUT <= x"000002120";
		when x"004aa" => DOUT <= x"000202141";
		when x"004ab" => DOUT <= x"000202140";
		when x"004ac" => DOUT <= x"000003121";
		when x"004ad" => DOUT <= x"0000031a0";
		when x"004ae" => DOUT <= x"0002031c1";
		when x"004af" => DOUT <= x"0002031c0";
		when x"004b0" => DOUT <= x"0000021a1";
		when x"004b1" => DOUT <= x"000002120";
		when x"004b2" => DOUT <= x"000202141";
		when x"004b3" => DOUT <= x"000202140";
		when x"004b4" => DOUT <= x"000003121";
		when x"004b5" => DOUT <= x"0000031a0";
		when x"004b6" => DOUT <= x"0002031c1";
		when x"004b7" => DOUT <= x"0002031c0";
		when x"004b8" => DOUT <= x"0000021a1";
		when x"004b9" => DOUT <= x"000002120";
		when x"004ba" => DOUT <= x"000202141";
		when x"004bb" => DOUT <= x"000202140";
		when x"004bc" => DOUT <= x"000003121";
		when x"004bd" => DOUT <= x"0000031a0";
		when x"004be" => DOUT <= x"0002031c1";
		when x"004bf" => DOUT <= x"0002031c0";
		when x"004c0" => DOUT <= x"0000021a1";
		when x"004c1" => DOUT <= x"000002120";
		when x"004c2" => DOUT <= x"000202141";
		when x"004c3" => DOUT <= x"000202140";
		when x"004c4" => DOUT <= x"000003121";
		when x"004c5" => DOUT <= x"0000031a0";
		when x"004c6" => DOUT <= x"0002031c1";
		when x"004c7" => DOUT <= x"0002031c0";
		when x"004c8" => DOUT <= x"0000021a1";
		when x"004c9" => DOUT <= x"000002120";
		when x"004ca" => DOUT <= x"000202141";
		when x"004cb" => DOUT <= x"000202140";
		when x"004cc" => DOUT <= x"000003121";
		when x"004cd" => DOUT <= x"0000031a0";
		when x"004ce" => DOUT <= x"0002031c1";
		when x"004cf" => DOUT <= x"0002031c0";
		when x"004d0" => DOUT <= x"0000021a1";
		when x"004d1" => DOUT <= x"000002120";
		when x"004d2" => DOUT <= x"000202141";
		when x"004d3" => DOUT <= x"000202140";
		when x"004d4" => DOUT <= x"000003121";
		when x"004d5" => DOUT <= x"0000031a0";
		when x"004d6" => DOUT <= x"0002031c1";
		when x"004d7" => DOUT <= x"0002031c0";
		when x"004d8" => DOUT <= x"0000021a1";
		when x"004d9" => DOUT <= x"000002120";
		when x"004da" => DOUT <= x"000202141";
		when x"004db" => DOUT <= x"000202140";
		when x"004dc" => DOUT <= x"000003121";
		when x"004dd" => DOUT <= x"0000031a0";
		when x"004de" => DOUT <= x"0002031c1";
		when x"004df" => DOUT <= x"0002031c0";
		when x"004e0" => DOUT <= x"0000021a1";
		when x"004e1" => DOUT <= x"000002120";
		when x"004e2" => DOUT <= x"000202141";
		when x"004e3" => DOUT <= x"000202140";
		when x"004e4" => DOUT <= x"000003121";
		when x"004e5" => DOUT <= x"0000031a0";
		when x"004e6" => DOUT <= x"0002031c1";
		when x"004e7" => DOUT <= x"0002031c0";
		when x"004e8" => DOUT <= x"0000021a1";
		when x"004e9" => DOUT <= x"000002120";
		when x"004ea" => DOUT <= x"000202141";
		when x"004eb" => DOUT <= x"000202140";
		when x"004ec" => DOUT <= x"000003121";
		when x"004ed" => DOUT <= x"0000031a0";
		when x"004ee" => DOUT <= x"0002031c1";
		when x"004ef" => DOUT <= x"0002031c0";
		when x"004f0" => DOUT <= x"0000021a1";
		when x"004f1" => DOUT <= x"000002120";
		when x"004f2" => DOUT <= x"000202141";
		when x"004f3" => DOUT <= x"000202140";
		when x"004f4" => DOUT <= x"000003121";
		when x"004f5" => DOUT <= x"0000031a0";
		when x"004f6" => DOUT <= x"0002031c1";
		when x"004f7" => DOUT <= x"0002031c0";
		when x"004f8" => DOUT <= x"0000021a1";
		when x"004f9" => DOUT <= x"000002120";
		when x"004fa" => DOUT <= x"000202141";
		when x"004fb" => DOUT <= x"000202140";
		when x"004fc" => DOUT <= x"000003121";
		when x"004fd" => DOUT <= x"0000031a0";
		when x"004fe" => DOUT <= x"0002031c1";
		when x"004ff" => DOUT <= x"0002031c0";
		when x"00500" => DOUT <= x"0000021a1";
		when x"00501" => DOUT <= x"000002120";
		when x"00502" => DOUT <= x"000202141";
		when x"00503" => DOUT <= x"000202140";
		when x"00504" => DOUT <= x"000003121";
		when x"00505" => DOUT <= x"0000031a0";
		when x"00506" => DOUT <= x"0002031c1";
		when x"00507" => DOUT <= x"0002031c0";
		when x"00508" => DOUT <= x"0000021a1";
		when x"00509" => DOUT <= x"000002120";
		when x"0050a" => DOUT <= x"000202141";
		when x"0050b" => DOUT <= x"000202140";
		when x"0050c" => DOUT <= x"000003121";
		when x"0050d" => DOUT <= x"0000031a0";
		when x"0050e" => DOUT <= x"0002031c1";
		when x"0050f" => DOUT <= x"0002031c0";
		when x"00510" => DOUT <= x"0000021a1";
		when x"00511" => DOUT <= x"000002120";
		when x"00512" => DOUT <= x"000202141";
		when x"00513" => DOUT <= x"000202140";
		when x"00514" => DOUT <= x"000003121";
		when x"00515" => DOUT <= x"0000031a0";
		when x"00516" => DOUT <= x"0002031c1";
		when x"00517" => DOUT <= x"0002031c0";
		when x"00518" => DOUT <= x"0000021a1";
		when x"00519" => DOUT <= x"000002120";
		when x"0051a" => DOUT <= x"000202141";
		when x"0051b" => DOUT <= x"000202140";
		when x"0051c" => DOUT <= x"000003121";
		when x"0051d" => DOUT <= x"0000031a0";
		when x"0051e" => DOUT <= x"0002031c1";
		when x"0051f" => DOUT <= x"0002031c0";
		when x"00520" => DOUT <= x"0000021a1";
		when x"00521" => DOUT <= x"000002120";
		when x"00522" => DOUT <= x"000202141";
		when x"00523" => DOUT <= x"000202140";
		when x"00524" => DOUT <= x"000003121";
		when x"00525" => DOUT <= x"0000031a0";
		when x"00526" => DOUT <= x"0002031c1";
		when x"00527" => DOUT <= x"0002031c0";
		when x"00528" => DOUT <= x"0000021a1";
		when x"00529" => DOUT <= x"000002120";
		when x"0052a" => DOUT <= x"000202141";
		when x"0052b" => DOUT <= x"000202140";
		when x"0052c" => DOUT <= x"000003121";
		when x"0052d" => DOUT <= x"0000031a0";
		when x"0052e" => DOUT <= x"0002031c1";
		when x"0052f" => DOUT <= x"0002031c0";
		when x"00530" => DOUT <= x"0000021a1";
		when x"00531" => DOUT <= x"000002120";
		when x"00532" => DOUT <= x"000202141";
		when x"00533" => DOUT <= x"000202140";
		when x"00534" => DOUT <= x"000003121";
		when x"00535" => DOUT <= x"0000031a0";
		when x"00536" => DOUT <= x"0002031c1";
		when x"00537" => DOUT <= x"0002031c0";
		when x"00538" => DOUT <= x"0000021a1";
		when x"00539" => DOUT <= x"000002120";
		when x"0053a" => DOUT <= x"000202141";
		when x"0053b" => DOUT <= x"000202140";
		when x"0053c" => DOUT <= x"000003121";
		when x"0053d" => DOUT <= x"0000031a0";
		when x"0053e" => DOUT <= x"0002031c1";
		when x"0053f" => DOUT <= x"0002031c0";
		when x"00540" => DOUT <= x"0000021a1";
		when x"00541" => DOUT <= x"000002120";
		when x"00542" => DOUT <= x"000202141";
		when x"00543" => DOUT <= x"000202140";
		when x"00544" => DOUT <= x"000003121";
		when x"00545" => DOUT <= x"0000031a0";
		when x"00546" => DOUT <= x"0002031c1";
		when x"00547" => DOUT <= x"0002031c0";
		when x"00548" => DOUT <= x"0000021a1";
		when x"00549" => DOUT <= x"000002120";
		when x"0054a" => DOUT <= x"000202141";
		when x"0054b" => DOUT <= x"000202140";
		when x"0054c" => DOUT <= x"000003121";
		when x"0054d" => DOUT <= x"0000031a0";
		when x"0054e" => DOUT <= x"0002031c1";
		when x"0054f" => DOUT <= x"0002031c0";
		when x"00550" => DOUT <= x"0000021a1";
		when x"00551" => DOUT <= x"000002120";
		when x"00552" => DOUT <= x"000202141";
		when x"00553" => DOUT <= x"000202140";
		when x"00554" => DOUT <= x"000003121";
		when x"00555" => DOUT <= x"0000031a0";
		when x"00556" => DOUT <= x"0002031c1";
		when x"00557" => DOUT <= x"0002031c0";
		when x"00558" => DOUT <= x"0000021a1";
		when x"00559" => DOUT <= x"000002120";
		when x"0055a" => DOUT <= x"000202141";
		when x"0055b" => DOUT <= x"000202140";
		when x"0055c" => DOUT <= x"000003121";
		when x"0055d" => DOUT <= x"0000031a0";
		when x"0055e" => DOUT <= x"0002031c1";
		when x"0055f" => DOUT <= x"0002031c0";
		when x"00560" => DOUT <= x"0000021a1";
		when x"00561" => DOUT <= x"000002120";
		when x"00562" => DOUT <= x"000202141";
		when x"00563" => DOUT <= x"000202140";
		when x"00564" => DOUT <= x"000003121";
		when x"00565" => DOUT <= x"0000031a0";
		when x"00566" => DOUT <= x"0002031c1";
		when x"00567" => DOUT <= x"0002031c0";
		when x"00568" => DOUT <= x"0000021a1";
		when x"00569" => DOUT <= x"000002120";
		when x"0056a" => DOUT <= x"000202141";
		when x"0056b" => DOUT <= x"000202140";
		when x"0056c" => DOUT <= x"000003121";
		when x"0056d" => DOUT <= x"0000031a0";
		when x"0056e" => DOUT <= x"0002031c1";
		when x"0056f" => DOUT <= x"0002031c0";
		when x"00570" => DOUT <= x"0000021a1";
		when x"00571" => DOUT <= x"000002120";
		when x"00572" => DOUT <= x"000202141";
		when x"00573" => DOUT <= x"000202140";
		when x"00574" => DOUT <= x"000003121";
		when x"00575" => DOUT <= x"0000031a0";
		when x"00576" => DOUT <= x"0002031c1";
		when x"00577" => DOUT <= x"0002031c0";
		when x"00578" => DOUT <= x"0000021a1";
		when x"00579" => DOUT <= x"000002120";
		when x"0057a" => DOUT <= x"000202141";
		when x"0057b" => DOUT <= x"000202140";
		when x"0057c" => DOUT <= x"000003121";
		when x"0057d" => DOUT <= x"0000031a0";
		when x"0057e" => DOUT <= x"0002031c1";
		when x"0057f" => DOUT <= x"0002031c0";
		when x"00580" => DOUT <= x"0000021a1";
		when x"00581" => DOUT <= x"000002120";
		when x"00582" => DOUT <= x"000202141";
		when x"00583" => DOUT <= x"000202140";
		when x"00584" => DOUT <= x"000003121";
		when x"00585" => DOUT <= x"0000031a0";
		when x"00586" => DOUT <= x"0002031c1";
		when x"00587" => DOUT <= x"0002031c0";
		when x"00588" => DOUT <= x"0000021a1";
		when x"00589" => DOUT <= x"000002120";
		when x"0058a" => DOUT <= x"000202141";
		when x"0058b" => DOUT <= x"000202140";
		when x"0058c" => DOUT <= x"000003121";
		when x"0058d" => DOUT <= x"0000031a0";
		when x"0058e" => DOUT <= x"0002031c1";
		when x"0058f" => DOUT <= x"0002031c0";
		when x"00590" => DOUT <= x"0000021a1";
		when x"00591" => DOUT <= x"000002120";
		when x"00592" => DOUT <= x"000202141";
		when x"00593" => DOUT <= x"000202140";
		when x"00594" => DOUT <= x"000003121";
		when x"00595" => DOUT <= x"0000031a0";
		when x"00596" => DOUT <= x"0002031c1";
		when x"00597" => DOUT <= x"0002031c0";
		when x"00598" => DOUT <= x"0000021a1";
		when x"00599" => DOUT <= x"000002120";
		when x"0059a" => DOUT <= x"000202141";
		when x"0059b" => DOUT <= x"000202140";
		when x"0059c" => DOUT <= x"000003121";
		when x"0059d" => DOUT <= x"0000031a0";
		when x"0059e" => DOUT <= x"0002031c1";
		when x"0059f" => DOUT <= x"0002031c0";
		when x"005a0" => DOUT <= x"0000021a1";
		when x"005a1" => DOUT <= x"000002120";
		when x"005a2" => DOUT <= x"000202141";
		when x"005a3" => DOUT <= x"000202140";
		when x"005a4" => DOUT <= x"000003121";
		when x"005a5" => DOUT <= x"0000031a0";
		when x"005a6" => DOUT <= x"0002031c1";
		when x"005a7" => DOUT <= x"0002031c0";
		when x"005a8" => DOUT <= x"0000021a1";
		when x"005a9" => DOUT <= x"000002120";
		when x"005aa" => DOUT <= x"000202141";
		when x"005ab" => DOUT <= x"000202140";
		when x"005ac" => DOUT <= x"000003121";
		when x"005ad" => DOUT <= x"0000031a0";
		when x"005ae" => DOUT <= x"0002031c1";
		when x"005af" => DOUT <= x"0002031c0";
		when x"005b0" => DOUT <= x"0000021a1";
		when x"005b1" => DOUT <= x"000002120";
		when x"005b2" => DOUT <= x"000202141";
		when x"005b3" => DOUT <= x"000202140";
		when x"005b4" => DOUT <= x"000003121";
		when x"005b5" => DOUT <= x"0000031a0";
		when x"005b6" => DOUT <= x"0002031c1";
		when x"005b7" => DOUT <= x"0002031c0";
		when x"005b8" => DOUT <= x"0000021a1";
		when x"005b9" => DOUT <= x"000002120";
		when x"005ba" => DOUT <= x"000202141";
		when x"005bb" => DOUT <= x"000202140";
		when x"005bc" => DOUT <= x"000003121";
		when x"005bd" => DOUT <= x"0000031a0";
		when x"005be" => DOUT <= x"0002031c1";
		when x"005bf" => DOUT <= x"0002031c0";
		when x"005c0" => DOUT <= x"0000021a1";
		when x"005c1" => DOUT <= x"000002120";
		when x"005c2" => DOUT <= x"000202141";
		when x"005c3" => DOUT <= x"000202140";
		when x"005c4" => DOUT <= x"000003121";
		when x"005c5" => DOUT <= x"0000031a0";
		when x"005c6" => DOUT <= x"0002031c1";
		when x"005c7" => DOUT <= x"0002031c0";
		when x"005c8" => DOUT <= x"0000021a1";
		when x"005c9" => DOUT <= x"000002120";
		when x"005ca" => DOUT <= x"000202141";
		when x"005cb" => DOUT <= x"000202140";
		when x"005cc" => DOUT <= x"000003121";
		when x"005cd" => DOUT <= x"0000031a0";
		when x"005ce" => DOUT <= x"0002031c1";
		when x"005cf" => DOUT <= x"0002031c0";
		when x"005d0" => DOUT <= x"0000021a1";
		when x"005d1" => DOUT <= x"000002120";
		when x"005d2" => DOUT <= x"000202141";
		when x"005d3" => DOUT <= x"000202140";
		when x"005d4" => DOUT <= x"000003121";
		when x"005d5" => DOUT <= x"0000031a0";
		when x"005d6" => DOUT <= x"0002031c1";
		when x"005d7" => DOUT <= x"0002031c0";
		when x"005d8" => DOUT <= x"0000021a1";
		when x"005d9" => DOUT <= x"000002120";
		when x"005da" => DOUT <= x"000202141";
		when x"005db" => DOUT <= x"000202140";
		when x"005dc" => DOUT <= x"000003121";
		when x"005dd" => DOUT <= x"0000031a0";
		when x"005de" => DOUT <= x"0002031c1";
		when x"005df" => DOUT <= x"0002031c0";
		when x"005e0" => DOUT <= x"0000021a1";
		when x"005e1" => DOUT <= x"000002120";
		when x"005e2" => DOUT <= x"000202141";
		when x"005e3" => DOUT <= x"000202140";
		when x"005e4" => DOUT <= x"000003121";
		when x"005e5" => DOUT <= x"0000031a0";
		when x"005e6" => DOUT <= x"0002031c1";
		when x"005e7" => DOUT <= x"0002031c0";
		when x"005e8" => DOUT <= x"0000021a1";
		when x"005e9" => DOUT <= x"000002120";
		when x"005ea" => DOUT <= x"000202141";
		when x"005eb" => DOUT <= x"000202140";
		when x"005ec" => DOUT <= x"000003121";
		when x"005ed" => DOUT <= x"0000031a0";
		when x"005ee" => DOUT <= x"0002031c1";
		when x"005ef" => DOUT <= x"0002031c0";
		when x"005f0" => DOUT <= x"0000021a1";
		when x"005f1" => DOUT <= x"000002120";
		when x"005f2" => DOUT <= x"000202141";
		when x"005f3" => DOUT <= x"000202140";
		when x"005f4" => DOUT <= x"000003121";
		when x"005f5" => DOUT <= x"0000031a0";
		when x"005f6" => DOUT <= x"0002031c1";
		when x"005f7" => DOUT <= x"0002031c0";
		when x"005f8" => DOUT <= x"0000021a1";
		when x"005f9" => DOUT <= x"000002120";
		when x"005fa" => DOUT <= x"000202141";
		when x"005fb" => DOUT <= x"000202140";
		when x"005fc" => DOUT <= x"000003121";
		when x"005fd" => DOUT <= x"0000031a0";
		when x"005fe" => DOUT <= x"0002031c1";
		when x"005ff" => DOUT <= x"0002031c0";
		when x"00600" => DOUT <= x"0000021a1";
		when x"00601" => DOUT <= x"000002120";
		when x"00602" => DOUT <= x"000202141";
		when x"00603" => DOUT <= x"000202140";
		when x"00604" => DOUT <= x"000003121";
		when x"00605" => DOUT <= x"0000031a0";
		when x"00606" => DOUT <= x"0002031c1";
		when x"00607" => DOUT <= x"0002031c0";
		when x"00608" => DOUT <= x"0000021a1";
		when x"00609" => DOUT <= x"000002120";
		when x"0060a" => DOUT <= x"000202141";
		when x"0060b" => DOUT <= x"000202140";
		when x"0060c" => DOUT <= x"000003121";
		when x"0060d" => DOUT <= x"0000031a0";
		when x"0060e" => DOUT <= x"0002031c1";
		when x"0060f" => DOUT <= x"0002031c0";
		when x"00610" => DOUT <= x"0000021a1";
		when x"00611" => DOUT <= x"000002120";
		when x"00612" => DOUT <= x"000202141";
		when x"00613" => DOUT <= x"000202140";
		when x"00614" => DOUT <= x"000003121";
		when x"00615" => DOUT <= x"0000031a0";
		when x"00616" => DOUT <= x"0002031c1";
		when x"00617" => DOUT <= x"0002031c0";
		when x"00618" => DOUT <= x"0000021a1";
		when x"00619" => DOUT <= x"000002120";
		when x"0061a" => DOUT <= x"000202141";
		when x"0061b" => DOUT <= x"000202140";
		when x"0061c" => DOUT <= x"000003121";
		when x"0061d" => DOUT <= x"0000031a0";
		when x"0061e" => DOUT <= x"0002031c1";
		when x"0061f" => DOUT <= x"0002031c0";
		when x"00620" => DOUT <= x"0000021a1";
		when x"00621" => DOUT <= x"000002120";
		when x"00622" => DOUT <= x"000202141";
		when x"00623" => DOUT <= x"000202140";
		when x"00624" => DOUT <= x"000003121";
		when x"00625" => DOUT <= x"0000031a0";
		when x"00626" => DOUT <= x"0002031c1";
		when x"00627" => DOUT <= x"0002031c0";
		when x"00628" => DOUT <= x"0000021a1";
		when x"00629" => DOUT <= x"000002120";
		when x"0062a" => DOUT <= x"000202141";
		when x"0062b" => DOUT <= x"000202140";
		when x"0062c" => DOUT <= x"000003121";
		when x"0062d" => DOUT <= x"0000031a0";
		when x"0062e" => DOUT <= x"0002031c1";
		when x"0062f" => DOUT <= x"0002031c0";
		when x"00630" => DOUT <= x"0000021a1";
		when x"00631" => DOUT <= x"000002120";
		when x"00632" => DOUT <= x"000202141";
		when x"00633" => DOUT <= x"000202140";
		when x"00634" => DOUT <= x"000003121";
		when x"00635" => DOUT <= x"0000031a0";
		when x"00636" => DOUT <= x"0002031c1";
		when x"00637" => DOUT <= x"0002031c0";
		when x"00638" => DOUT <= x"0000021a1";
		when x"00639" => DOUT <= x"000002120";
		when x"0063a" => DOUT <= x"000202141";
		when x"0063b" => DOUT <= x"000202140";
		when x"0063c" => DOUT <= x"000003121";
		when x"0063d" => DOUT <= x"0000031a0";
		when x"0063e" => DOUT <= x"0002031c1";
		when x"0063f" => DOUT <= x"0002031c0";
		when x"00640" => DOUT <= x"0000021a1";
		when x"00641" => DOUT <= x"000002120";
		when x"00642" => DOUT <= x"000202141";
		when x"00643" => DOUT <= x"000202140";
		when x"00644" => DOUT <= x"000003121";
		when x"00645" => DOUT <= x"0000031a0";
		when x"00646" => DOUT <= x"0002031c1";
		when x"00647" => DOUT <= x"0002031c0";
		when x"00648" => DOUT <= x"0000021a1";
		when x"00649" => DOUT <= x"000002120";
		when x"0064a" => DOUT <= x"000202141";
		when x"0064b" => DOUT <= x"000202140";
		when x"0064c" => DOUT <= x"000003121";
		when x"0064d" => DOUT <= x"0000031a0";
		when x"0064e" => DOUT <= x"0002031c1";
		when x"0064f" => DOUT <= x"0002031c0";
		when x"00650" => DOUT <= x"0000021a1";
		when x"00651" => DOUT <= x"000002120";
		when x"00652" => DOUT <= x"000202141";
		when x"00653" => DOUT <= x"000202140";
		when x"00654" => DOUT <= x"000003121";
		when x"00655" => DOUT <= x"0000031a0";
		when x"00656" => DOUT <= x"0002031c1";
		when x"00657" => DOUT <= x"0002031c0";
		when x"00658" => DOUT <= x"0000021a1";
		when x"00659" => DOUT <= x"000002120";
		when x"0065a" => DOUT <= x"000202141";
		when x"0065b" => DOUT <= x"000202140";
		when x"0065c" => DOUT <= x"000003121";
		when x"0065d" => DOUT <= x"0000031a0";
		when x"0065e" => DOUT <= x"0002031c1";
		when x"0065f" => DOUT <= x"0002031c0";
		when x"00660" => DOUT <= x"0000021a1";
		when x"00661" => DOUT <= x"000002120";
		when x"00662" => DOUT <= x"000202141";
		when x"00663" => DOUT <= x"000202140";
		when x"00664" => DOUT <= x"000003121";
		when x"00665" => DOUT <= x"0000031a0";
		when x"00666" => DOUT <= x"0002031c1";
		when x"00667" => DOUT <= x"0002031c0";
		when x"00668" => DOUT <= x"0000021a1";
		when x"00669" => DOUT <= x"000002120";
		when x"0066a" => DOUT <= x"000202141";
		when x"0066b" => DOUT <= x"000202140";
		when x"0066c" => DOUT <= x"000003121";
		when x"0066d" => DOUT <= x"0000031a0";
		when x"0066e" => DOUT <= x"0002031c1";
		when x"0066f" => DOUT <= x"0002031c0";
		when x"00670" => DOUT <= x"0000021a1";
		when x"00671" => DOUT <= x"000002120";
		when x"00672" => DOUT <= x"000202141";
		when x"00673" => DOUT <= x"000202140";
		when x"00674" => DOUT <= x"000003121";
		when x"00675" => DOUT <= x"0000031a0";
		when x"00676" => DOUT <= x"0002031c1";
		when x"00677" => DOUT <= x"0002031c0";
		when x"00678" => DOUT <= x"0000021a1";
		when x"00679" => DOUT <= x"000002120";
		when x"0067a" => DOUT <= x"000202141";
		when x"0067b" => DOUT <= x"000202140";
		when x"0067c" => DOUT <= x"000003121";
		when x"0067d" => DOUT <= x"0000031a0";
		when x"0067e" => DOUT <= x"0002031c1";
		when x"0067f" => DOUT <= x"0002031c0";
		when x"00680" => DOUT <= x"0000021a1";
		when x"00681" => DOUT <= x"000002120";
		when x"00682" => DOUT <= x"000202141";
		when x"00683" => DOUT <= x"000202140";
		when x"00684" => DOUT <= x"000003121";
		when x"00685" => DOUT <= x"0000031a0";
		when x"00686" => DOUT <= x"0002031c1";
		when x"00687" => DOUT <= x"0002031c0";
		when x"00688" => DOUT <= x"0000021a1";
		when x"00689" => DOUT <= x"000002120";
		when x"0068a" => DOUT <= x"000202141";
		when x"0068b" => DOUT <= x"000202140";
		when x"0068c" => DOUT <= x"000003121";
		when x"0068d" => DOUT <= x"0000031a0";
		when x"0068e" => DOUT <= x"0002031c1";
		when x"0068f" => DOUT <= x"0002031c0";
		when x"00690" => DOUT <= x"0000021a1";
		when x"00691" => DOUT <= x"000002120";
		when x"00692" => DOUT <= x"000202141";
		when x"00693" => DOUT <= x"000202140";
		when x"00694" => DOUT <= x"000003121";
		when x"00695" => DOUT <= x"0000031a0";
		when x"00696" => DOUT <= x"0002031c1";
		when x"00697" => DOUT <= x"0002031c0";
		when x"00698" => DOUT <= x"0000021a1";
		when x"00699" => DOUT <= x"000002120";
		when x"0069a" => DOUT <= x"000202141";
		when x"0069b" => DOUT <= x"000202140";
		when x"0069c" => DOUT <= x"000003121";
		when x"0069d" => DOUT <= x"0000031a0";
		when x"0069e" => DOUT <= x"0002031c1";
		when x"0069f" => DOUT <= x"0002031c0";
		when x"006a0" => DOUT <= x"0000021a1";
		when x"006a1" => DOUT <= x"000002120";
		when x"006a2" => DOUT <= x"000202141";
		when x"006a3" => DOUT <= x"000202140";
		when x"006a4" => DOUT <= x"000003121";
		when x"006a5" => DOUT <= x"0000031a0";
		when x"006a6" => DOUT <= x"0002031c1";
		when x"006a7" => DOUT <= x"0002031c0";
		when x"006a8" => DOUT <= x"0000021a1";
		when x"006a9" => DOUT <= x"000002120";
		when x"006aa" => DOUT <= x"000202141";
		when x"006ab" => DOUT <= x"000202140";
		when x"006ac" => DOUT <= x"000003121";
		when x"006ad" => DOUT <= x"0000031a0";
		when x"006ae" => DOUT <= x"0002031c1";
		when x"006af" => DOUT <= x"0002031c0";
		when x"006b0" => DOUT <= x"0000021a1";
		when x"006b1" => DOUT <= x"000002120";
		when x"006b2" => DOUT <= x"000202141";
		when x"006b3" => DOUT <= x"000202140";
		when x"006b4" => DOUT <= x"000003121";
		when x"006b5" => DOUT <= x"0000031a0";
		when x"006b6" => DOUT <= x"0002031c1";
		when x"006b7" => DOUT <= x"0002031c0";
		when x"006b8" => DOUT <= x"0000021a1";
		when x"006b9" => DOUT <= x"000002120";
		when x"006ba" => DOUT <= x"000202141";
		when x"006bb" => DOUT <= x"000202140";
		when x"006bc" => DOUT <= x"000003121";
		when x"006bd" => DOUT <= x"0000031a0";
		when x"006be" => DOUT <= x"0002031c1";
		when x"006bf" => DOUT <= x"0002031c0";
		when x"006c0" => DOUT <= x"0000021a1";
		when x"006c1" => DOUT <= x"000002120";
		when x"006c2" => DOUT <= x"000202141";
		when x"006c3" => DOUT <= x"000202140";
		when x"006c4" => DOUT <= x"000003121";
		when x"006c5" => DOUT <= x"0000031a0";
		when x"006c6" => DOUT <= x"0002031c1";
		when x"006c7" => DOUT <= x"0002031c0";
		when x"006c8" => DOUT <= x"0000021a1";
		when x"006c9" => DOUT <= x"000002120";
		when x"006ca" => DOUT <= x"000202141";
		when x"006cb" => DOUT <= x"000202140";
		when x"006cc" => DOUT <= x"000003121";
		when x"006cd" => DOUT <= x"0000031a0";
		when x"006ce" => DOUT <= x"0002031c1";
		when x"006cf" => DOUT <= x"0002031c0";
		when x"006d0" => DOUT <= x"0000021a1";
		when x"006d1" => DOUT <= x"000002120";
		when x"006d2" => DOUT <= x"000202141";
		when x"006d3" => DOUT <= x"000202140";
		when x"006d4" => DOUT <= x"000003121";
		when x"006d5" => DOUT <= x"0000031a0";
		when x"006d6" => DOUT <= x"0002031c1";
		when x"006d7" => DOUT <= x"0002031c0";
		when x"006d8" => DOUT <= x"0000021a1";
		when x"006d9" => DOUT <= x"000002120";
		when x"006da" => DOUT <= x"000202141";
		when x"006db" => DOUT <= x"000202140";
		when x"006dc" => DOUT <= x"000003121";
		when x"006dd" => DOUT <= x"0000031a0";
		when x"006de" => DOUT <= x"0002031c1";
		when x"006df" => DOUT <= x"0002031c0";
		when x"006e0" => DOUT <= x"0000021a1";
		when x"006e1" => DOUT <= x"000002120";
		when x"006e2" => DOUT <= x"000202141";
		when x"006e3" => DOUT <= x"000202140";
		when x"006e4" => DOUT <= x"000003121";
		when x"006e5" => DOUT <= x"0000031a0";
		when x"006e6" => DOUT <= x"0002031c1";
		when x"006e7" => DOUT <= x"0002031c0";
		when x"006e8" => DOUT <= x"0000021a1";
		when x"006e9" => DOUT <= x"000002120";
		when x"006ea" => DOUT <= x"000202141";
		when x"006eb" => DOUT <= x"000202140";
		when x"006ec" => DOUT <= x"000003121";
		when x"006ed" => DOUT <= x"0000031a0";
		when x"006ee" => DOUT <= x"0002031c1";
		when x"006ef" => DOUT <= x"0002031c0";
		when x"006f0" => DOUT <= x"0000021a1";
		when x"006f1" => DOUT <= x"000002120";
		when x"006f2" => DOUT <= x"000202141";
		when x"006f3" => DOUT <= x"000202140";
		when x"006f4" => DOUT <= x"000003121";
		when x"006f5" => DOUT <= x"0000031a0";
		when x"006f6" => DOUT <= x"0002031c1";
		when x"006f7" => DOUT <= x"0002031c0";
		when x"006f8" => DOUT <= x"0000021a1";
		when x"006f9" => DOUT <= x"000002120";
		when x"006fa" => DOUT <= x"000202141";
		when x"006fb" => DOUT <= x"000202140";
		when x"006fc" => DOUT <= x"000003121";
		when x"006fd" => DOUT <= x"0000031a0";
		when x"006fe" => DOUT <= x"0002031c1";
		when x"006ff" => DOUT <= x"0002031c0";
		when x"00700" => DOUT <= x"0000021a1";
		when x"00701" => DOUT <= x"000002120";
		when x"00702" => DOUT <= x"000202141";
		when x"00703" => DOUT <= x"000202140";
		when x"00704" => DOUT <= x"000003121";
		when x"00705" => DOUT <= x"0000031a0";
		when x"00706" => DOUT <= x"0002031c1";
		when x"00707" => DOUT <= x"0002031c0";
		when x"00708" => DOUT <= x"0000021a1";
		when x"00709" => DOUT <= x"000002120";
		when x"0070a" => DOUT <= x"000202141";
		when x"0070b" => DOUT <= x"000202140";
		when x"0070c" => DOUT <= x"000003121";
		when x"0070d" => DOUT <= x"0000031a0";
		when x"0070e" => DOUT <= x"0002031c1";
		when x"0070f" => DOUT <= x"0002031c0";
		when x"00710" => DOUT <= x"0000021a1";
		when x"00711" => DOUT <= x"000002120";
		when x"00712" => DOUT <= x"000202141";
		when x"00713" => DOUT <= x"000202140";
		when x"00714" => DOUT <= x"000003121";
		when x"00715" => DOUT <= x"0000031a0";
		when x"00716" => DOUT <= x"0002031c1";
		when x"00717" => DOUT <= x"0002031c0";
		when x"00718" => DOUT <= x"0000021a1";
		when x"00719" => DOUT <= x"000002120";
		when x"0071a" => DOUT <= x"000202141";
		when x"0071b" => DOUT <= x"000202140";
		when x"0071c" => DOUT <= x"000003121";
		when x"0071d" => DOUT <= x"0000031a0";
		when x"0071e" => DOUT <= x"0002031c1";
		when x"0071f" => DOUT <= x"0002031c0";
		when x"00720" => DOUT <= x"0000021a1";
		when x"00721" => DOUT <= x"000002120";
		when x"00722" => DOUT <= x"000202141";
		when x"00723" => DOUT <= x"000202140";
		when x"00724" => DOUT <= x"000003121";
		when x"00725" => DOUT <= x"0000031a0";
		when x"00726" => DOUT <= x"0002031c1";
		when x"00727" => DOUT <= x"0002031c0";
		when x"00728" => DOUT <= x"0000021a1";
		when x"00729" => DOUT <= x"000002120";
		when x"0072a" => DOUT <= x"000202141";
		when x"0072b" => DOUT <= x"000202140";
		when x"0072c" => DOUT <= x"000003121";
		when x"0072d" => DOUT <= x"0000031a0";
		when x"0072e" => DOUT <= x"0002031c1";
		when x"0072f" => DOUT <= x"0002031c0";
		when x"00730" => DOUT <= x"0000021a1";
		when x"00731" => DOUT <= x"000002120";
		when x"00732" => DOUT <= x"000202141";
		when x"00733" => DOUT <= x"000202140";
		when x"00734" => DOUT <= x"000003121";
		when x"00735" => DOUT <= x"0000031a0";
		when x"00736" => DOUT <= x"0002031c1";
		when x"00737" => DOUT <= x"0002031c0";
		when x"00738" => DOUT <= x"0000021a1";
		when x"00739" => DOUT <= x"000002120";
		when x"0073a" => DOUT <= x"000202141";
		when x"0073b" => DOUT <= x"000202140";
		when x"0073c" => DOUT <= x"000003121";
		when x"0073d" => DOUT <= x"0000031a0";
		when x"0073e" => DOUT <= x"0002031c1";
		when x"0073f" => DOUT <= x"0002031c0";
		when x"00740" => DOUT <= x"0000021a1";
		when x"00741" => DOUT <= x"000002120";
		when x"00742" => DOUT <= x"000202141";
		when x"00743" => DOUT <= x"000202140";
		when x"00744" => DOUT <= x"000003121";
		when x"00745" => DOUT <= x"0000031a0";
		when x"00746" => DOUT <= x"0002031c1";
		when x"00747" => DOUT <= x"0002031c0";
		when x"00748" => DOUT <= x"0000021a1";
		when x"00749" => DOUT <= x"000002120";
		when x"0074a" => DOUT <= x"000202141";
		when x"0074b" => DOUT <= x"000202140";
		when x"0074c" => DOUT <= x"000003121";
		when x"0074d" => DOUT <= x"0000031a0";
		when x"0074e" => DOUT <= x"0002031c1";
		when x"0074f" => DOUT <= x"0002031c0";
		when x"00750" => DOUT <= x"0000021a1";
		when x"00751" => DOUT <= x"000002120";
		when x"00752" => DOUT <= x"000202141";
		when x"00753" => DOUT <= x"000202140";
		when x"00754" => DOUT <= x"000003121";
		when x"00755" => DOUT <= x"0000031a0";
		when x"00756" => DOUT <= x"0002031c1";
		when x"00757" => DOUT <= x"0002031c0";
		when x"00758" => DOUT <= x"0000021a1";
		when x"00759" => DOUT <= x"000002120";
		when x"0075a" => DOUT <= x"000202141";
		when x"0075b" => DOUT <= x"000202140";
		when x"0075c" => DOUT <= x"000003121";
		when x"0075d" => DOUT <= x"0000031a0";
		when x"0075e" => DOUT <= x"0002031c1";
		when x"0075f" => DOUT <= x"0002031c0";
		when x"00760" => DOUT <= x"0000021a1";
		when x"00761" => DOUT <= x"000002120";
		when x"00762" => DOUT <= x"000202141";
		when x"00763" => DOUT <= x"000202140";
		when x"00764" => DOUT <= x"000003121";
		when x"00765" => DOUT <= x"0000031a0";
		when x"00766" => DOUT <= x"0002031c1";
		when x"00767" => DOUT <= x"0002031c0";
		when x"00768" => DOUT <= x"0000021a1";
		when x"00769" => DOUT <= x"000002120";
		when x"0076a" => DOUT <= x"000202141";
		when x"0076b" => DOUT <= x"000202140";
		when x"0076c" => DOUT <= x"000003121";
		when x"0076d" => DOUT <= x"0000031a0";
		when x"0076e" => DOUT <= x"0002031c1";
		when x"0076f" => DOUT <= x"0002031c0";
		when x"00770" => DOUT <= x"0000021a1";
		when x"00771" => DOUT <= x"000002120";
		when x"00772" => DOUT <= x"000202141";
		when x"00773" => DOUT <= x"000202140";
		when x"00774" => DOUT <= x"000003121";
		when x"00775" => DOUT <= x"0000031a0";
		when x"00776" => DOUT <= x"0002031c1";
		when x"00777" => DOUT <= x"0002031c0";
		when x"00778" => DOUT <= x"0000021a1";
		when x"00779" => DOUT <= x"000002120";
		when x"0077a" => DOUT <= x"000202141";
		when x"0077b" => DOUT <= x"000202140";
		when x"0077c" => DOUT <= x"000003121";
		when x"0077d" => DOUT <= x"0000031a0";
		when x"0077e" => DOUT <= x"0002031c1";
		when x"0077f" => DOUT <= x"0002031c0";
		when x"00780" => DOUT <= x"0000021a1";
		when x"00781" => DOUT <= x"000002120";
		when x"00782" => DOUT <= x"000202141";
		when x"00783" => DOUT <= x"000202140";
		when x"00784" => DOUT <= x"000003121";
		when x"00785" => DOUT <= x"0000031a0";
		when x"00786" => DOUT <= x"0002031c1";
		when x"00787" => DOUT <= x"0002031c0";
		when x"00788" => DOUT <= x"0000021a1";
		when x"00789" => DOUT <= x"000002120";
		when x"0078a" => DOUT <= x"000202141";
		when x"0078b" => DOUT <= x"000202140";
		when x"0078c" => DOUT <= x"000003121";
		when x"0078d" => DOUT <= x"0000031a0";
		when x"0078e" => DOUT <= x"0002031c1";
		when x"0078f" => DOUT <= x"0002031c0";
		when x"00790" => DOUT <= x"0000021a1";
		when x"00791" => DOUT <= x"000002120";
		when x"00792" => DOUT <= x"000202141";
		when x"00793" => DOUT <= x"000202140";
		when x"00794" => DOUT <= x"000003121";
		when x"00795" => DOUT <= x"0000031a0";
		when x"00796" => DOUT <= x"0002031c1";
		when x"00797" => DOUT <= x"0002031c0";
		when x"00798" => DOUT <= x"0000021a1";
		when x"00799" => DOUT <= x"000002120";
		when x"0079a" => DOUT <= x"000202141";
		when x"0079b" => DOUT <= x"000202140";
		when x"0079c" => DOUT <= x"000003121";
		when x"0079d" => DOUT <= x"0000031a0";
		when x"0079e" => DOUT <= x"0002031c1";
		when x"0079f" => DOUT <= x"0002031c0";
		when x"007a0" => DOUT <= x"0000021a1";
		when x"007a1" => DOUT <= x"000002120";
		when x"007a2" => DOUT <= x"000202141";
		when x"007a3" => DOUT <= x"000202140";
		when x"007a4" => DOUT <= x"000003121";
		when x"007a5" => DOUT <= x"0000031a0";
		when x"007a6" => DOUT <= x"0002031c1";
		when x"007a7" => DOUT <= x"0002031c0";
		when x"007a8" => DOUT <= x"0000021a1";
		when x"007a9" => DOUT <= x"000002120";
		when x"007aa" => DOUT <= x"000202141";
		when x"007ab" => DOUT <= x"000202140";
		when x"007ac" => DOUT <= x"000003121";
		when x"007ad" => DOUT <= x"0000031a0";
		when x"007ae" => DOUT <= x"0002031c1";
		when x"007af" => DOUT <= x"0002031c0";
		when x"007b0" => DOUT <= x"0000021a1";
		when x"007b1" => DOUT <= x"000002120";
		when x"007b2" => DOUT <= x"000202141";
		when x"007b3" => DOUT <= x"000202140";
		when x"007b4" => DOUT <= x"000003121";
		when x"007b5" => DOUT <= x"0000031a0";
		when x"007b6" => DOUT <= x"0002031c1";
		when x"007b7" => DOUT <= x"0002031c0";
		when x"007b8" => DOUT <= x"0000021a1";
		when x"007b9" => DOUT <= x"000002120";
		when x"007ba" => DOUT <= x"000202141";
		when x"007bb" => DOUT <= x"000202140";
		when x"007bc" => DOUT <= x"000003121";
		when x"007bd" => DOUT <= x"0000031a0";
		when x"007be" => DOUT <= x"0002031c1";
		when x"007bf" => DOUT <= x"0002031c0";
		when x"007c0" => DOUT <= x"0000021a1";
		when x"007c1" => DOUT <= x"000002120";
		when x"007c2" => DOUT <= x"000202141";
		when x"007c3" => DOUT <= x"000202140";
		when x"007c4" => DOUT <= x"000003121";
		when x"007c5" => DOUT <= x"0000031a0";
		when x"007c6" => DOUT <= x"0002031c1";
		when x"007c7" => DOUT <= x"0002031c0";
		when x"007c8" => DOUT <= x"0000021a1";
		when x"007c9" => DOUT <= x"000002120";
		when x"007ca" => DOUT <= x"000202141";
		when x"007cb" => DOUT <= x"000202140";
		when x"007cc" => DOUT <= x"000003121";
		when x"007cd" => DOUT <= x"0000031a0";
		when x"007ce" => DOUT <= x"0002031c1";
		when x"007cf" => DOUT <= x"0002031c0";
		when x"007d0" => DOUT <= x"0000021a1";
		when x"007d1" => DOUT <= x"000002120";
		when x"007d2" => DOUT <= x"000202141";
		when x"007d3" => DOUT <= x"000202140";
		when x"007d4" => DOUT <= x"000003121";
		when x"007d5" => DOUT <= x"0000031a0";
		when x"007d6" => DOUT <= x"0002031c1";
		when x"007d7" => DOUT <= x"0002031c0";
		when x"007d8" => DOUT <= x"0000021a1";
		when x"007d9" => DOUT <= x"000002120";
		when x"007da" => DOUT <= x"000202141";
		when x"007db" => DOUT <= x"000202140";
		when x"007dc" => DOUT <= x"000003121";
		when x"007dd" => DOUT <= x"0000031a0";
		when x"007de" => DOUT <= x"0002031c1";
		when x"007df" => DOUT <= x"0002031c0";
		when x"007e0" => DOUT <= x"0000021a1";
		when x"007e1" => DOUT <= x"000002120";
		when x"007e2" => DOUT <= x"000202141";
		when x"007e3" => DOUT <= x"000202140";
		when x"007e4" => DOUT <= x"000003121";
		when x"007e5" => DOUT <= x"0000031a0";
		when x"007e6" => DOUT <= x"0002031c1";
		when x"007e7" => DOUT <= x"0002031c0";
		when x"007e8" => DOUT <= x"0000021a1";
		when x"007e9" => DOUT <= x"000002120";
		when x"007ea" => DOUT <= x"000202141";
		when x"007eb" => DOUT <= x"000202140";
		when x"007ec" => DOUT <= x"000003121";
		when x"007ed" => DOUT <= x"0000031a0";
		when x"007ee" => DOUT <= x"0002031c1";
		when x"007ef" => DOUT <= x"0002031c0";
		when x"007f0" => DOUT <= x"0000021a1";
		when x"007f1" => DOUT <= x"000002120";
		when x"007f2" => DOUT <= x"000202141";
		when x"007f3" => DOUT <= x"000202140";
		when x"007f4" => DOUT <= x"000003121";
		when x"007f5" => DOUT <= x"0000031a0";
		when x"007f6" => DOUT <= x"0002031c1";
		when x"007f7" => DOUT <= x"0002031c0";
		when x"007f8" => DOUT <= x"0000021a1";
		when x"007f9" => DOUT <= x"000002120";
		when x"007fa" => DOUT <= x"000202141";
		when x"007fb" => DOUT <= x"000202140";
		when x"007fc" => DOUT <= x"000003121";
		when x"007fd" => DOUT <= x"0000031a0";
		when x"007fe" => DOUT <= x"0002031c1";
		when x"007ff" => DOUT <= x"0002031c0";
		when x"00800" => DOUT <= x"0000021a1";
		when x"00801" => DOUT <= x"000002120";
		when x"00802" => DOUT <= x"000202141";
		when x"00803" => DOUT <= x"000202140";
		when x"00804" => DOUT <= x"000003121";
		when x"00805" => DOUT <= x"0000031a0";
		when x"00806" => DOUT <= x"0002031c1";
		when x"00807" => DOUT <= x"0002031c0";
		when x"00808" => DOUT <= x"0000021a1";
		when x"00809" => DOUT <= x"000002120";
		when x"0080a" => DOUT <= x"000202141";
		when x"0080b" => DOUT <= x"000202140";
		when x"0080c" => DOUT <= x"000003121";
		when x"0080d" => DOUT <= x"0000031a0";
		when x"0080e" => DOUT <= x"0002031c1";
		when x"0080f" => DOUT <= x"0002031c0";
		when x"00810" => DOUT <= x"0000021a1";
		when x"00811" => DOUT <= x"000002120";
		when x"00812" => DOUT <= x"000202141";
		when x"00813" => DOUT <= x"000202140";
		when x"00814" => DOUT <= x"000003121";
		when x"00815" => DOUT <= x"0000031a0";
		when x"00816" => DOUT <= x"0002031c1";
		when x"00817" => DOUT <= x"0002031c0";
		when x"00818" => DOUT <= x"0000021a1";
		when x"00819" => DOUT <= x"000002120";
		when x"0081a" => DOUT <= x"000202141";
		when x"0081b" => DOUT <= x"000202140";
		when x"0081c" => DOUT <= x"000003121";
		when x"0081d" => DOUT <= x"0000031a0";
		when x"0081e" => DOUT <= x"0002031c1";
		when x"0081f" => DOUT <= x"0002031c0";
		when x"00820" => DOUT <= x"0000021a1";
		when x"00821" => DOUT <= x"000002120";
		when x"00822" => DOUT <= x"000202141";
		when x"00823" => DOUT <= x"000202140";
		when x"00824" => DOUT <= x"000003121";
		when x"00825" => DOUT <= x"0000031a0";
		when x"00826" => DOUT <= x"0002031c1";
		when x"00827" => DOUT <= x"0002031c0";
		when x"00828" => DOUT <= x"0000021a1";
		when x"00829" => DOUT <= x"000002120";
		when x"0082a" => DOUT <= x"000202141";
		when x"0082b" => DOUT <= x"000202140";
		when x"0082c" => DOUT <= x"000003121";
		when x"0082d" => DOUT <= x"0000031a0";
		when x"0082e" => DOUT <= x"0002031c1";
		when x"0082f" => DOUT <= x"0002031c0";
		when x"00830" => DOUT <= x"0000021a1";
		when x"00831" => DOUT <= x"000002120";
		when x"00832" => DOUT <= x"000202141";
		when x"00833" => DOUT <= x"000202140";
		when x"00834" => DOUT <= x"000003121";
		when x"00835" => DOUT <= x"0000031a0";
		when x"00836" => DOUT <= x"0002031c1";
		when x"00837" => DOUT <= x"0002031c0";
		when x"00838" => DOUT <= x"0000021a1";
		when x"00839" => DOUT <= x"000002120";
		when x"0083a" => DOUT <= x"000202141";
		when x"0083b" => DOUT <= x"000202140";
		when x"0083c" => DOUT <= x"000003121";
		when x"0083d" => DOUT <= x"0000031a0";
		when x"0083e" => DOUT <= x"0002031c1";
		when x"0083f" => DOUT <= x"0002031c0";
		when x"00840" => DOUT <= x"0000021a1";
		when x"00841" => DOUT <= x"000002120";
		when x"00842" => DOUT <= x"000202141";
		when x"00843" => DOUT <= x"000202140";
		when x"00844" => DOUT <= x"000003121";
		when x"00845" => DOUT <= x"0000031a0";
		when x"00846" => DOUT <= x"0002031c1";
		when x"00847" => DOUT <= x"0002031c0";
		when x"00848" => DOUT <= x"0000021a1";
		when x"00849" => DOUT <= x"000002120";
		when x"0084a" => DOUT <= x"000202141";
		when x"0084b" => DOUT <= x"000202140";
		when x"0084c" => DOUT <= x"000003121";
		when x"0084d" => DOUT <= x"0000031a0";
		when x"0084e" => DOUT <= x"0002031c1";
		when x"0084f" => DOUT <= x"0002031c0";
		when x"00850" => DOUT <= x"0000021a1";
		when x"00851" => DOUT <= x"000002120";
		when x"00852" => DOUT <= x"000202141";
		when x"00853" => DOUT <= x"000202140";
		when x"00854" => DOUT <= x"000003121";
		when x"00855" => DOUT <= x"0000031a0";
		when x"00856" => DOUT <= x"0002031c1";
		when x"00857" => DOUT <= x"0002031c0";
		when x"00858" => DOUT <= x"0000021a1";
		when x"00859" => DOUT <= x"000002120";
		when x"0085a" => DOUT <= x"000202141";
		when x"0085b" => DOUT <= x"000202140";
		when x"0085c" => DOUT <= x"000003121";
		when x"0085d" => DOUT <= x"0000031a0";
		when x"0085e" => DOUT <= x"0002031c1";
		when x"0085f" => DOUT <= x"0002031c0";
		when x"00860" => DOUT <= x"0000021a1";
		when x"00861" => DOUT <= x"000002120";
		when x"00862" => DOUT <= x"000202141";
		when x"00863" => DOUT <= x"000202140";
		when x"00864" => DOUT <= x"000003121";
		when x"00865" => DOUT <= x"0000031a0";
		when x"00866" => DOUT <= x"0002031c1";
		when x"00867" => DOUT <= x"0002031c0";
		when x"00868" => DOUT <= x"0000021a1";
		when x"00869" => DOUT <= x"000002120";
		when x"0086a" => DOUT <= x"000202141";
		when x"0086b" => DOUT <= x"000202140";
		when x"0086c" => DOUT <= x"000003121";
		when x"0086d" => DOUT <= x"0000031a0";
		when x"0086e" => DOUT <= x"0002031c1";
		when x"0086f" => DOUT <= x"0002031c0";
		when x"00870" => DOUT <= x"0000021a1";
		when x"00871" => DOUT <= x"000002120";
		when x"00872" => DOUT <= x"000202141";
		when x"00873" => DOUT <= x"000202140";
		when x"00874" => DOUT <= x"000003121";
		when x"00875" => DOUT <= x"0000031a0";
		when x"00876" => DOUT <= x"0002031c1";
		when x"00877" => DOUT <= x"0002031c0";
		when x"00878" => DOUT <= x"0000021a1";
		when x"00879" => DOUT <= x"000002120";
		when x"0087a" => DOUT <= x"000202141";
		when x"0087b" => DOUT <= x"000202140";
		when x"0087c" => DOUT <= x"000003121";
		when x"0087d" => DOUT <= x"0000031a0";
		when x"0087e" => DOUT <= x"0002031c1";
		when x"0087f" => DOUT <= x"0002031c0";
		when x"00880" => DOUT <= x"0000021a1";
		when x"00881" => DOUT <= x"000002120";
		when x"00882" => DOUT <= x"000202141";
		when x"00883" => DOUT <= x"000202140";
		when x"00884" => DOUT <= x"000003121";
		when x"00885" => DOUT <= x"0000031a0";
		when x"00886" => DOUT <= x"0002031c1";
		when x"00887" => DOUT <= x"0002031c0";
		when x"00888" => DOUT <= x"0000021a1";
		when x"00889" => DOUT <= x"000002120";
		when x"0088a" => DOUT <= x"000202141";
		when x"0088b" => DOUT <= x"000202140";
		when x"0088c" => DOUT <= x"000003121";
		when x"0088d" => DOUT <= x"0000031a0";
		when x"0088e" => DOUT <= x"0002031c1";
		when x"0088f" => DOUT <= x"0002031c0";
		when x"00890" => DOUT <= x"0000021a1";
		when x"00891" => DOUT <= x"000002120";
		when x"00892" => DOUT <= x"000202141";
		when x"00893" => DOUT <= x"000202140";
		when x"00894" => DOUT <= x"000003121";
		when x"00895" => DOUT <= x"0000031a0";
		when x"00896" => DOUT <= x"0002031c1";
		when x"00897" => DOUT <= x"0002031c0";
		when x"00898" => DOUT <= x"0000021a1";
		when x"00899" => DOUT <= x"000002120";
		when x"0089a" => DOUT <= x"000202141";
		when x"0089b" => DOUT <= x"000202140";
		when x"0089c" => DOUT <= x"000003121";
		when x"0089d" => DOUT <= x"0000031a0";
		when x"0089e" => DOUT <= x"0002031c1";
		when x"0089f" => DOUT <= x"0002031c0";
		when x"008a0" => DOUT <= x"0000021a1";
		when x"008a1" => DOUT <= x"000002120";
		when x"008a2" => DOUT <= x"000202141";
		when x"008a3" => DOUT <= x"000202140";
		when x"008a4" => DOUT <= x"000003121";
		when x"008a5" => DOUT <= x"0000031a0";
		when x"008a6" => DOUT <= x"0002031c1";
		when x"008a7" => DOUT <= x"0002031c0";
		when x"008a8" => DOUT <= x"0000021a1";
		when x"008a9" => DOUT <= x"000002120";
		when x"008aa" => DOUT <= x"000202141";
		when x"008ab" => DOUT <= x"000202140";
		when x"008ac" => DOUT <= x"000003121";
		when x"008ad" => DOUT <= x"0000031a0";
		when x"008ae" => DOUT <= x"0002031c1";
		when x"008af" => DOUT <= x"0002031c0";
		when x"008b0" => DOUT <= x"0000021a1";
		when x"008b1" => DOUT <= x"000002120";
		when x"008b2" => DOUT <= x"000202141";
		when x"008b3" => DOUT <= x"000202140";
		when x"008b4" => DOUT <= x"000003121";
		when x"008b5" => DOUT <= x"0000031a0";
		when x"008b6" => DOUT <= x"0002031c1";
		when x"008b7" => DOUT <= x"0002031c0";
		when x"008b8" => DOUT <= x"0000021a1";
		when x"008b9" => DOUT <= x"000002120";
		when x"008ba" => DOUT <= x"000202141";
		when x"008bb" => DOUT <= x"000202140";
		when x"008bc" => DOUT <= x"000003121";
		when x"008bd" => DOUT <= x"0000031a0";
		when x"008be" => DOUT <= x"0002031c1";
		when x"008bf" => DOUT <= x"0002031c0";
		when x"008c0" => DOUT <= x"0000021a1";
		when x"008c1" => DOUT <= x"000002120";
		when x"008c2" => DOUT <= x"000202141";
		when x"008c3" => DOUT <= x"000202140";
		when x"008c4" => DOUT <= x"000003121";
		when x"008c5" => DOUT <= x"0000031a0";
		when x"008c6" => DOUT <= x"0002031c1";
		when x"008c7" => DOUT <= x"0002031c0";
		when x"008c8" => DOUT <= x"0000021a1";
		when x"008c9" => DOUT <= x"000002120";
		when x"008ca" => DOUT <= x"000202141";
		when x"008cb" => DOUT <= x"000202140";
		when x"008cc" => DOUT <= x"000003121";
		when x"008cd" => DOUT <= x"0000031a0";
		when x"008ce" => DOUT <= x"0002031c1";
		when x"008cf" => DOUT <= x"0002031c0";
		when x"008d0" => DOUT <= x"0000021a1";
		when x"008d1" => DOUT <= x"000002120";
		when x"008d2" => DOUT <= x"000202141";
		when x"008d3" => DOUT <= x"000202140";
		when x"008d4" => DOUT <= x"000003121";
		when x"008d5" => DOUT <= x"0000031a0";
		when x"008d6" => DOUT <= x"0002031c1";
		when x"008d7" => DOUT <= x"0002031c0";
		when x"008d8" => DOUT <= x"0000021a1";
		when x"008d9" => DOUT <= x"000002120";
		when x"008da" => DOUT <= x"000202141";
		when x"008db" => DOUT <= x"000202140";
		when x"008dc" => DOUT <= x"000003121";
		when x"008dd" => DOUT <= x"0000031a0";
		when x"008de" => DOUT <= x"0002031c1";
		when x"008df" => DOUT <= x"0002031c0";
		when x"008e0" => DOUT <= x"0000021a1";
		when x"008e1" => DOUT <= x"000002120";
		when x"008e2" => DOUT <= x"000202141";
		when x"008e3" => DOUT <= x"000202140";
		when x"008e4" => DOUT <= x"000003121";
		when x"008e5" => DOUT <= x"0000031a0";
		when x"008e6" => DOUT <= x"0002031c1";
		when x"008e7" => DOUT <= x"0002031c0";
		when x"008e8" => DOUT <= x"0000021a1";
		when x"008e9" => DOUT <= x"000002120";
		when x"008ea" => DOUT <= x"000202141";
		when x"008eb" => DOUT <= x"000202140";
		when x"008ec" => DOUT <= x"000003121";
		when x"008ed" => DOUT <= x"0000031a0";
		when x"008ee" => DOUT <= x"0002031c1";
		when x"008ef" => DOUT <= x"0002031c0";
		when x"008f0" => DOUT <= x"0000021a1";
		when x"008f1" => DOUT <= x"000002120";
		when x"008f2" => DOUT <= x"000202141";
		when x"008f3" => DOUT <= x"000202140";
		when x"008f4" => DOUT <= x"000003121";
		when x"008f5" => DOUT <= x"0000031a0";
		when x"008f6" => DOUT <= x"0002031c1";
		when x"008f7" => DOUT <= x"0002031c0";
		when x"008f8" => DOUT <= x"0000021a1";
		when x"008f9" => DOUT <= x"000002120";
		when x"008fa" => DOUT <= x"000202141";
		when x"008fb" => DOUT <= x"000202140";
		when x"008fc" => DOUT <= x"000003121";
		when x"008fd" => DOUT <= x"0000031a0";
		when x"008fe" => DOUT <= x"0002031c1";
		when x"008ff" => DOUT <= x"0002031c0";
		when x"00900" => DOUT <= x"0000021a1";
		when x"00901" => DOUT <= x"000002120";
		when x"00902" => DOUT <= x"000202141";
		when x"00903" => DOUT <= x"000202140";
		when x"00904" => DOUT <= x"000003121";
		when x"00905" => DOUT <= x"0000031a0";
		when x"00906" => DOUT <= x"0002031c1";
		when x"00907" => DOUT <= x"0002031c0";
		when x"00908" => DOUT <= x"0000021a1";
		when x"00909" => DOUT <= x"000002120";
		when x"0090a" => DOUT <= x"000202141";
		when x"0090b" => DOUT <= x"000202140";
		when x"0090c" => DOUT <= x"000003121";
		when x"0090d" => DOUT <= x"0000031a0";
		when x"0090e" => DOUT <= x"0002031c1";
		when x"0090f" => DOUT <= x"0002031c0";
		when x"00910" => DOUT <= x"0000021a1";
		when x"00911" => DOUT <= x"000002120";
		when x"00912" => DOUT <= x"000202141";
		when x"00913" => DOUT <= x"000202140";
		when x"00914" => DOUT <= x"000003121";
		when x"00915" => DOUT <= x"0000031a0";
		when x"00916" => DOUT <= x"0002031c1";
		when x"00917" => DOUT <= x"0002031c0";
		when x"00918" => DOUT <= x"0000021a1";
		when x"00919" => DOUT <= x"000002120";
		when x"0091a" => DOUT <= x"000202141";
		when x"0091b" => DOUT <= x"000202140";
		when x"0091c" => DOUT <= x"000003121";
		when x"0091d" => DOUT <= x"0000031a0";
		when x"0091e" => DOUT <= x"0002031c1";
		when x"0091f" => DOUT <= x"0002031c0";
		when x"00920" => DOUT <= x"0000021a1";
		when x"00921" => DOUT <= x"000002120";
		when x"00922" => DOUT <= x"000202141";
		when x"00923" => DOUT <= x"000202140";
		when x"00924" => DOUT <= x"000003121";
		when x"00925" => DOUT <= x"0000031a0";
		when x"00926" => DOUT <= x"0002031c1";
		when x"00927" => DOUT <= x"0002031c0";
		when x"00928" => DOUT <= x"0000021a1";
		when x"00929" => DOUT <= x"000002120";
		when x"0092a" => DOUT <= x"000202141";
		when x"0092b" => DOUT <= x"000202140";
		when x"0092c" => DOUT <= x"000003121";
		when x"0092d" => DOUT <= x"0000031a0";
		when x"0092e" => DOUT <= x"0002031c1";
		when x"0092f" => DOUT <= x"0002031c0";
		when x"00930" => DOUT <= x"0000021a1";
		when x"00931" => DOUT <= x"000002120";
		when x"00932" => DOUT <= x"000202141";
		when x"00933" => DOUT <= x"000202140";
		when x"00934" => DOUT <= x"000003121";
		when x"00935" => DOUT <= x"0000031a0";
		when x"00936" => DOUT <= x"0002031c1";
		when x"00937" => DOUT <= x"0002031c0";
		when x"00938" => DOUT <= x"0000021a1";
		when x"00939" => DOUT <= x"000002120";
		when x"0093a" => DOUT <= x"000202141";
		when x"0093b" => DOUT <= x"000202140";
		when x"0093c" => DOUT <= x"000003121";
		when x"0093d" => DOUT <= x"0000031a0";
		when x"0093e" => DOUT <= x"0002031c1";
		when x"0093f" => DOUT <= x"0002031c0";
		when x"00940" => DOUT <= x"0000021a1";
		when x"00941" => DOUT <= x"000002120";
		when x"00942" => DOUT <= x"000202141";
		when x"00943" => DOUT <= x"000202140";
		when x"00944" => DOUT <= x"000003121";
		when x"00945" => DOUT <= x"0000031a0";
		when x"00946" => DOUT <= x"0002031c1";
		when x"00947" => DOUT <= x"0002031c0";
		when x"00948" => DOUT <= x"0000021a1";
		when x"00949" => DOUT <= x"000002120";
		when x"0094a" => DOUT <= x"000202141";
		when x"0094b" => DOUT <= x"000202140";
		when x"0094c" => DOUT <= x"000003121";
		when x"0094d" => DOUT <= x"0000031a0";
		when x"0094e" => DOUT <= x"0002031c1";
		when x"0094f" => DOUT <= x"0002031c0";
		when x"00950" => DOUT <= x"0000021a1";
		when x"00951" => DOUT <= x"000002120";
		when x"00952" => DOUT <= x"000202141";
		when x"00953" => DOUT <= x"000202140";
		when x"00954" => DOUT <= x"000003121";
		when x"00955" => DOUT <= x"0000031a0";
		when x"00956" => DOUT <= x"0002031c1";
		when x"00957" => DOUT <= x"0002031c0";
		when x"00958" => DOUT <= x"0000021a1";
		when x"00959" => DOUT <= x"000002120";
		when x"0095a" => DOUT <= x"000202141";
		when x"0095b" => DOUT <= x"000202140";
		when x"0095c" => DOUT <= x"000003121";
		when x"0095d" => DOUT <= x"0000031a0";
		when x"0095e" => DOUT <= x"0002031c1";
		when x"0095f" => DOUT <= x"0002031c0";
		when x"00960" => DOUT <= x"0000021a1";
		when x"00961" => DOUT <= x"000002120";
		when x"00962" => DOUT <= x"000202141";
		when x"00963" => DOUT <= x"000202140";
		when x"00964" => DOUT <= x"000003121";
		when x"00965" => DOUT <= x"0000031a0";
		when x"00966" => DOUT <= x"0002031c1";
		when x"00967" => DOUT <= x"0002031c0";
		when x"00968" => DOUT <= x"0000021a1";
		when x"00969" => DOUT <= x"000002120";
		when x"0096a" => DOUT <= x"000202141";
		when x"0096b" => DOUT <= x"000202140";
		when x"0096c" => DOUT <= x"000003121";
		when x"0096d" => DOUT <= x"0000031a0";
		when x"0096e" => DOUT <= x"0002031c1";
		when x"0096f" => DOUT <= x"0002031c0";
		when x"00970" => DOUT <= x"0000021a1";
		when x"00971" => DOUT <= x"000002120";
		when x"00972" => DOUT <= x"000202141";
		when x"00973" => DOUT <= x"000202140";
		when x"00974" => DOUT <= x"000003121";
		when x"00975" => DOUT <= x"0000031a0";
		when x"00976" => DOUT <= x"0002031c1";
		when x"00977" => DOUT <= x"0002031c0";
		when x"00978" => DOUT <= x"0000021a1";
		when x"00979" => DOUT <= x"000002120";
		when x"0097a" => DOUT <= x"000202141";
		when x"0097b" => DOUT <= x"000202140";
		when x"0097c" => DOUT <= x"000003121";
		when x"0097d" => DOUT <= x"0000031a0";
		when x"0097e" => DOUT <= x"0002031c1";
		when x"0097f" => DOUT <= x"0002031c0";
		when x"00980" => DOUT <= x"0000021a1";
		when x"00981" => DOUT <= x"000002120";
		when x"00982" => DOUT <= x"000202141";
		when x"00983" => DOUT <= x"000202140";
		when x"00984" => DOUT <= x"000003121";
		when x"00985" => DOUT <= x"0000031a0";
		when x"00986" => DOUT <= x"0002031c1";
		when x"00987" => DOUT <= x"0002031c0";
		when x"00988" => DOUT <= x"0000021a1";
		when x"00989" => DOUT <= x"000002120";
		when x"0098a" => DOUT <= x"000202141";
		when x"0098b" => DOUT <= x"000202140";
		when x"0098c" => DOUT <= x"000003121";
		when x"0098d" => DOUT <= x"0000031a0";
		when x"0098e" => DOUT <= x"0002031c1";
		when x"0098f" => DOUT <= x"0002031c0";
		when x"00990" => DOUT <= x"0000021a1";
		when x"00991" => DOUT <= x"000002120";
		when x"00992" => DOUT <= x"000202141";
		when x"00993" => DOUT <= x"000202140";
		when x"00994" => DOUT <= x"000003121";
		when x"00995" => DOUT <= x"0000031a0";
		when x"00996" => DOUT <= x"0002031c1";
		when x"00997" => DOUT <= x"0002031c0";
		when x"00998" => DOUT <= x"0000021a1";
		when x"00999" => DOUT <= x"000002120";
		when x"0099a" => DOUT <= x"000202141";
		when x"0099b" => DOUT <= x"000202140";
		when x"0099c" => DOUT <= x"000003121";
		when x"0099d" => DOUT <= x"0000031a0";
		when x"0099e" => DOUT <= x"0002031c1";
		when x"0099f" => DOUT <= x"0002031c0";
		when x"009a0" => DOUT <= x"0000021a1";
		when x"009a1" => DOUT <= x"000002120";
		when x"009a2" => DOUT <= x"000202141";
		when x"009a3" => DOUT <= x"000202140";
		when x"009a4" => DOUT <= x"000003121";
		when x"009a5" => DOUT <= x"0000031a0";
		when x"009a6" => DOUT <= x"0002031c1";
		when x"009a7" => DOUT <= x"0002031c0";
		when x"009a8" => DOUT <= x"0000021a1";
		when x"009a9" => DOUT <= x"000002120";
		when x"009aa" => DOUT <= x"000202141";
		when x"009ab" => DOUT <= x"000202140";
		when x"009ac" => DOUT <= x"000003121";
		when x"009ad" => DOUT <= x"0000031a0";
		when x"009ae" => DOUT <= x"0002031c1";
		when x"009af" => DOUT <= x"0002031c0";
		when x"009b0" => DOUT <= x"0000021a1";
		when x"009b1" => DOUT <= x"000002120";
		when x"009b2" => DOUT <= x"000202141";
		when x"009b3" => DOUT <= x"000202140";
		when x"009b4" => DOUT <= x"000003121";
		when x"009b5" => DOUT <= x"0000031a0";
		when x"009b6" => DOUT <= x"0002031c1";
		when x"009b7" => DOUT <= x"0002031c0";
		when x"009b8" => DOUT <= x"0000021a1";
		when x"009b9" => DOUT <= x"000002120";
		when x"009ba" => DOUT <= x"000202141";
		when x"009bb" => DOUT <= x"000202140";
		when x"009bc" => DOUT <= x"000003121";
		when x"009bd" => DOUT <= x"0000031a0";
		when x"009be" => DOUT <= x"0002031c1";
		when x"009bf" => DOUT <= x"0002031c0";
		when x"009c0" => DOUT <= x"0000021a1";
		when x"009c1" => DOUT <= x"000002120";
		when x"009c2" => DOUT <= x"000202141";
		when x"009c3" => DOUT <= x"000202140";
		when x"009c4" => DOUT <= x"000003121";
		when x"009c5" => DOUT <= x"0000031a0";
		when x"009c6" => DOUT <= x"0002031c1";
		when x"009c7" => DOUT <= x"0002031c0";
		when x"009c8" => DOUT <= x"0000021a1";
		when x"009c9" => DOUT <= x"000002120";
		when x"009ca" => DOUT <= x"000202141";
		when x"009cb" => DOUT <= x"000202140";
		when x"009cc" => DOUT <= x"000003121";
		when x"009cd" => DOUT <= x"0000031a0";
		when x"009ce" => DOUT <= x"0002031c1";
		when x"009cf" => DOUT <= x"0002031c0";
		when x"009d0" => DOUT <= x"0000021a1";
		when x"009d1" => DOUT <= x"000002120";
		when x"009d2" => DOUT <= x"000202141";
		when x"009d3" => DOUT <= x"000202140";
		when x"009d4" => DOUT <= x"000003121";
		when x"009d5" => DOUT <= x"0000031a0";
		when x"009d6" => DOUT <= x"0002031c1";
		when x"009d7" => DOUT <= x"0002031c0";
		when x"009d8" => DOUT <= x"0000021a1";
		when x"009d9" => DOUT <= x"000002120";
		when x"009da" => DOUT <= x"000202141";
		when x"009db" => DOUT <= x"000202140";
		when x"009dc" => DOUT <= x"000003121";
		when x"009dd" => DOUT <= x"0000031a0";
		when x"009de" => DOUT <= x"0002031c1";
		when x"009df" => DOUT <= x"0002031c0";
		when x"009e0" => DOUT <= x"0000021a1";
		when x"009e1" => DOUT <= x"000002120";
		when x"009e2" => DOUT <= x"000202141";
		when x"009e3" => DOUT <= x"000202140";
		when x"009e4" => DOUT <= x"000003121";
		when x"009e5" => DOUT <= x"0000031a0";
		when x"009e6" => DOUT <= x"0002031c1";
		when x"009e7" => DOUT <= x"0002031c0";
		when x"009e8" => DOUT <= x"0000021a1";
		when x"009e9" => DOUT <= x"000002120";
		when x"009ea" => DOUT <= x"000202141";
		when x"009eb" => DOUT <= x"000202140";
		when x"009ec" => DOUT <= x"000003121";
		when x"009ed" => DOUT <= x"0000031a0";
		when x"009ee" => DOUT <= x"0002031c1";
		when x"009ef" => DOUT <= x"0002031c0";
		when x"009f0" => DOUT <= x"0000021a1";
		when x"009f1" => DOUT <= x"000002120";
		when x"009f2" => DOUT <= x"000202141";
		when x"009f3" => DOUT <= x"000202140";
		when x"009f4" => DOUT <= x"000003121";
		when x"009f5" => DOUT <= x"0000031a0";
		when x"009f6" => DOUT <= x"0002031c1";
		when x"009f7" => DOUT <= x"0002031c0";
		when x"009f8" => DOUT <= x"0000021a1";
		when x"009f9" => DOUT <= x"000002120";
		when x"009fa" => DOUT <= x"000202141";
		when x"009fb" => DOUT <= x"000202140";
		when x"009fc" => DOUT <= x"000003121";
		when x"009fd" => DOUT <= x"0000031a0";
		when x"009fe" => DOUT <= x"0002031c1";
		when x"009ff" => DOUT <= x"0002031c0";
		when x"00a00" => DOUT <= x"0000021a1";
		when x"00a01" => DOUT <= x"000002120";
		when x"00a02" => DOUT <= x"000202141";
		when x"00a03" => DOUT <= x"000202140";
		when x"00a04" => DOUT <= x"000003121";
		when x"00a05" => DOUT <= x"0000031a0";
		when x"00a06" => DOUT <= x"0002031c1";
		when x"00a07" => DOUT <= x"0002031c0";
		when x"00a08" => DOUT <= x"0000021a1";
		when x"00a09" => DOUT <= x"000002120";
		when x"00a0a" => DOUT <= x"000202141";
		when x"00a0b" => DOUT <= x"000202140";
		when x"00a0c" => DOUT <= x"000003121";
		when x"00a0d" => DOUT <= x"0000031a0";
		when x"00a0e" => DOUT <= x"0002031c1";
		when x"00a0f" => DOUT <= x"0002031c0";
		when x"00a10" => DOUT <= x"0000021a1";
		when x"00a11" => DOUT <= x"000002120";
		when x"00a12" => DOUT <= x"000202141";
		when x"00a13" => DOUT <= x"000202140";
		when x"00a14" => DOUT <= x"000003121";
		when x"00a15" => DOUT <= x"0000031a0";
		when x"00a16" => DOUT <= x"0002031c1";
		when x"00a17" => DOUT <= x"0002031c0";
		when x"00a18" => DOUT <= x"0000021a1";
		when x"00a19" => DOUT <= x"000002120";
		when x"00a1a" => DOUT <= x"000202141";
		when x"00a1b" => DOUT <= x"000202140";
		when x"00a1c" => DOUT <= x"000003121";
		when x"00a1d" => DOUT <= x"0000031a0";
		when x"00a1e" => DOUT <= x"0002031c1";
		when x"00a1f" => DOUT <= x"0002031c0";
		when x"00a20" => DOUT <= x"0000021a1";
		when x"00a21" => DOUT <= x"000002120";
		when x"00a22" => DOUT <= x"000202141";
		when x"00a23" => DOUT <= x"000202140";
		when x"00a24" => DOUT <= x"000003121";
		when x"00a25" => DOUT <= x"0000031a0";
		when x"00a26" => DOUT <= x"0002031c1";
		when x"00a27" => DOUT <= x"0002031c0";
		when x"00a28" => DOUT <= x"0000021a1";
		when x"00a29" => DOUT <= x"000002120";
		when x"00a2a" => DOUT <= x"000202141";
		when x"00a2b" => DOUT <= x"000202140";
		when x"00a2c" => DOUT <= x"000003121";
		when x"00a2d" => DOUT <= x"0000031a0";
		when x"00a2e" => DOUT <= x"0002031c1";
		when x"00a2f" => DOUT <= x"0002031c0";
		when x"00a30" => DOUT <= x"0000021a1";
		when x"00a31" => DOUT <= x"000002120";
		when x"00a32" => DOUT <= x"000202141";
		when x"00a33" => DOUT <= x"000202140";
		when x"00a34" => DOUT <= x"000003121";
		when x"00a35" => DOUT <= x"0000031a0";
		when x"00a36" => DOUT <= x"0002031c1";
		when x"00a37" => DOUT <= x"0002031c0";
		when x"00a38" => DOUT <= x"0000021a1";
		when x"00a39" => DOUT <= x"000002120";
		when x"00a3a" => DOUT <= x"000202141";
		when x"00a3b" => DOUT <= x"000202140";
		when x"00a3c" => DOUT <= x"000003121";
		when x"00a3d" => DOUT <= x"0000031a0";
		when x"00a3e" => DOUT <= x"0002031c1";
		when x"00a3f" => DOUT <= x"0002031c0";
		when x"00a40" => DOUT <= x"0000021a1";
		when x"00a41" => DOUT <= x"000002120";
		when x"00a42" => DOUT <= x"000202141";
		when x"00a43" => DOUT <= x"000202140";
		when x"00a44" => DOUT <= x"000003121";
		when x"00a45" => DOUT <= x"0000031a0";
		when x"00a46" => DOUT <= x"0002031c1";
		when x"00a47" => DOUT <= x"0002031c0";
		when x"00a48" => DOUT <= x"0000021a1";
		when x"00a49" => DOUT <= x"000002120";
		when x"00a4a" => DOUT <= x"000202141";
		when x"00a4b" => DOUT <= x"000202140";
		when x"00a4c" => DOUT <= x"000003121";
		when x"00a4d" => DOUT <= x"0000031a0";
		when x"00a4e" => DOUT <= x"0002031c1";
		when x"00a4f" => DOUT <= x"0002031c0";
		when x"00a50" => DOUT <= x"0000021a1";
		when x"00a51" => DOUT <= x"000002120";
		when x"00a52" => DOUT <= x"000202141";
		when x"00a53" => DOUT <= x"000202140";
		when x"00a54" => DOUT <= x"000003121";
		when x"00a55" => DOUT <= x"0000031a0";
		when x"00a56" => DOUT <= x"0002031c1";
		when x"00a57" => DOUT <= x"0002031c0";
		when x"00a58" => DOUT <= x"0000021a1";
		when x"00a59" => DOUT <= x"000002120";
		when x"00a5a" => DOUT <= x"000202141";
		when x"00a5b" => DOUT <= x"000202140";
		when x"00a5c" => DOUT <= x"000003121";
		when x"00a5d" => DOUT <= x"0000031a0";
		when x"00a5e" => DOUT <= x"0002031c1";
		when x"00a5f" => DOUT <= x"0002031c0";
		when x"00a60" => DOUT <= x"0000021a1";
		when x"00a61" => DOUT <= x"000002120";
		when x"00a62" => DOUT <= x"000202141";
		when x"00a63" => DOUT <= x"000202140";
		when x"00a64" => DOUT <= x"000003121";
		when x"00a65" => DOUT <= x"0000031a0";
		when x"00a66" => DOUT <= x"0002031c1";
		when x"00a67" => DOUT <= x"0002031c0";
		when x"00a68" => DOUT <= x"0000021a1";
		when x"00a69" => DOUT <= x"000002120";
		when x"00a6a" => DOUT <= x"000202141";
		when x"00a6b" => DOUT <= x"000202140";
		when x"00a6c" => DOUT <= x"000003121";
		when x"00a6d" => DOUT <= x"0000031a0";
		when x"00a6e" => DOUT <= x"0002031c1";
		when x"00a6f" => DOUT <= x"0002031c0";
		when x"00a70" => DOUT <= x"0000021a1";
		when x"00a71" => DOUT <= x"000002120";
		when x"00a72" => DOUT <= x"000202141";
		when x"00a73" => DOUT <= x"000202140";
		when x"00a74" => DOUT <= x"000003121";
		when x"00a75" => DOUT <= x"0000031a0";
		when x"00a76" => DOUT <= x"0002031c1";
		when x"00a77" => DOUT <= x"0002031c0";
		when x"00a78" => DOUT <= x"0000021a1";
		when x"00a79" => DOUT <= x"000002120";
		when x"00a7a" => DOUT <= x"000202141";
		when x"00a7b" => DOUT <= x"000202140";
		when x"00a7c" => DOUT <= x"000003121";
		when x"00a7d" => DOUT <= x"0000031a0";
		when x"00a7e" => DOUT <= x"0002031c1";
		when x"00a7f" => DOUT <= x"0002031c0";
		when x"00a80" => DOUT <= x"0000021a1";
		when x"00a81" => DOUT <= x"000002120";
		when x"00a82" => DOUT <= x"000202141";
		when x"00a83" => DOUT <= x"000202140";
		when x"00a84" => DOUT <= x"000003121";
		when x"00a85" => DOUT <= x"0000031a0";
		when x"00a86" => DOUT <= x"0002031c1";
		when x"00a87" => DOUT <= x"0002031c0";
		when x"00a88" => DOUT <= x"0000021a1";
		when x"00a89" => DOUT <= x"000002120";
		when x"00a8a" => DOUT <= x"000202141";
		when x"00a8b" => DOUT <= x"000202140";
		when x"00a8c" => DOUT <= x"000003121";
		when x"00a8d" => DOUT <= x"0000031a0";
		when x"00a8e" => DOUT <= x"0002031c1";
		when x"00a8f" => DOUT <= x"0002031c0";
		when x"00a90" => DOUT <= x"0000021a1";
		when x"00a91" => DOUT <= x"000002120";
		when x"00a92" => DOUT <= x"000202141";
		when x"00a93" => DOUT <= x"000202140";
		when x"00a94" => DOUT <= x"000003121";
		when x"00a95" => DOUT <= x"0000031a0";
		when x"00a96" => DOUT <= x"0002031c1";
		when x"00a97" => DOUT <= x"0002031c0";
		when x"00a98" => DOUT <= x"0000021a1";
		when x"00a99" => DOUT <= x"000002120";
		when x"00a9a" => DOUT <= x"000202141";
		when x"00a9b" => DOUT <= x"000202140";
		when x"00a9c" => DOUT <= x"000003121";
		when x"00a9d" => DOUT <= x"0000031a0";
		when x"00a9e" => DOUT <= x"0002031c1";
		when x"00a9f" => DOUT <= x"0002031c0";
		when x"00aa0" => DOUT <= x"0000021a1";
		when x"00aa1" => DOUT <= x"000002120";
		when x"00aa2" => DOUT <= x"000202141";
		when x"00aa3" => DOUT <= x"000202140";
		when x"00aa4" => DOUT <= x"000003121";
		when x"00aa5" => DOUT <= x"0000031a0";
		when x"00aa6" => DOUT <= x"0002031c1";
		when x"00aa7" => DOUT <= x"0002031c0";
		when x"00aa8" => DOUT <= x"0000021a1";
		when x"00aa9" => DOUT <= x"000002120";
		when x"00aaa" => DOUT <= x"000202141";
		when x"00aab" => DOUT <= x"000202140";
		when x"00aac" => DOUT <= x"000003121";
		when x"00aad" => DOUT <= x"0000031a0";
		when x"00aae" => DOUT <= x"0002031c1";
		when x"00aaf" => DOUT <= x"0002031c0";
		when x"00ab0" => DOUT <= x"0000021a1";
		when x"00ab1" => DOUT <= x"000002120";
		when x"00ab2" => DOUT <= x"000202141";
		when x"00ab3" => DOUT <= x"000202140";
		when x"00ab4" => DOUT <= x"000003121";
		when x"00ab5" => DOUT <= x"0000031a0";
		when x"00ab6" => DOUT <= x"0002031c1";
		when x"00ab7" => DOUT <= x"0002031c0";
		when x"00ab8" => DOUT <= x"0000021a1";
		when x"00ab9" => DOUT <= x"000002120";
		when x"00aba" => DOUT <= x"000202141";
		when x"00abb" => DOUT <= x"000202140";
		when x"00abc" => DOUT <= x"000003121";
		when x"00abd" => DOUT <= x"0000031a0";
		when x"00abe" => DOUT <= x"0002031c1";
		when x"00abf" => DOUT <= x"0002031c0";
		when x"00ac0" => DOUT <= x"0000021a1";
		when x"00ac1" => DOUT <= x"000002120";
		when x"00ac2" => DOUT <= x"000202141";
		when x"00ac3" => DOUT <= x"000202140";
		when x"00ac4" => DOUT <= x"000003121";
		when x"00ac5" => DOUT <= x"0000031a0";
		when x"00ac6" => DOUT <= x"0002031c1";
		when x"00ac7" => DOUT <= x"0002031c0";
		when x"00ac8" => DOUT <= x"0000021a1";
		when x"00ac9" => DOUT <= x"000002120";
		when x"00aca" => DOUT <= x"000202141";
		when x"00acb" => DOUT <= x"000202140";
		when x"00acc" => DOUT <= x"000003121";
		when x"00acd" => DOUT <= x"0000031a0";
		when x"00ace" => DOUT <= x"0002031c1";
		when x"00acf" => DOUT <= x"0002031c0";
		when x"00ad0" => DOUT <= x"0000021a1";
		when x"00ad1" => DOUT <= x"000002120";
		when x"00ad2" => DOUT <= x"000202141";
		when x"00ad3" => DOUT <= x"000202140";
		when x"00ad4" => DOUT <= x"000003121";
		when x"00ad5" => DOUT <= x"0000031a0";
		when x"00ad6" => DOUT <= x"0002031c1";
		when x"00ad7" => DOUT <= x"0002031c0";
		when x"00ad8" => DOUT <= x"0000021a1";
		when x"00ad9" => DOUT <= x"000002120";
		when x"00ada" => DOUT <= x"000202141";
		when x"00adb" => DOUT <= x"000202140";
		when x"00adc" => DOUT <= x"000003121";
		when x"00add" => DOUT <= x"0000031a0";
		when x"00ade" => DOUT <= x"0002031c1";
		when x"00adf" => DOUT <= x"0002031c0";
		when x"00ae0" => DOUT <= x"0000021a1";
		when x"00ae1" => DOUT <= x"000002120";
		when x"00ae2" => DOUT <= x"000202141";
		when x"00ae3" => DOUT <= x"000202140";
		when x"00ae4" => DOUT <= x"000003121";
		when x"00ae5" => DOUT <= x"0000031a0";
		when x"00ae6" => DOUT <= x"0002031c1";
		when x"00ae7" => DOUT <= x"0002031c0";
		when x"00ae8" => DOUT <= x"0000021a1";
		when x"00ae9" => DOUT <= x"000002120";
		when x"00aea" => DOUT <= x"000202141";
		when x"00aeb" => DOUT <= x"000202140";
		when x"00aec" => DOUT <= x"000003121";
		when x"00aed" => DOUT <= x"0000031a0";
		when x"00aee" => DOUT <= x"0002031c1";
		when x"00aef" => DOUT <= x"0002031c0";
		when x"00af0" => DOUT <= x"0000021a1";
		when x"00af1" => DOUT <= x"000002120";
		when x"00af2" => DOUT <= x"000202141";
		when x"00af3" => DOUT <= x"000202140";
		when x"00af4" => DOUT <= x"000003121";
		when x"00af5" => DOUT <= x"0000031a0";
		when x"00af6" => DOUT <= x"0002031c1";
		when x"00af7" => DOUT <= x"0002031c0";
		when x"00af8" => DOUT <= x"0000021a1";
		when x"00af9" => DOUT <= x"000002120";
		when x"00afa" => DOUT <= x"000202141";
		when x"00afb" => DOUT <= x"000202140";
		when x"00afc" => DOUT <= x"000003121";
		when x"00afd" => DOUT <= x"0000031a0";
		when x"00afe" => DOUT <= x"0002031c1";
		when x"00aff" => DOUT <= x"0002031c0";
		when x"00b00" => DOUT <= x"0000021a1";
		when x"00b01" => DOUT <= x"000002120";
		when x"00b02" => DOUT <= x"000202141";
		when x"00b03" => DOUT <= x"000202140";
		when x"00b04" => DOUT <= x"000003121";
		when x"00b05" => DOUT <= x"0000031a0";
		when x"00b06" => DOUT <= x"0002031c1";
		when x"00b07" => DOUT <= x"0002031c0";
		when x"00b08" => DOUT <= x"0000021a1";
		when x"00b09" => DOUT <= x"000002120";
		when x"00b0a" => DOUT <= x"000202141";
		when x"00b0b" => DOUT <= x"000202140";
		when x"00b0c" => DOUT <= x"000003121";
		when x"00b0d" => DOUT <= x"0000031a0";
		when x"00b0e" => DOUT <= x"0002031c1";
		when x"00b0f" => DOUT <= x"0002031c0";
		when x"00b10" => DOUT <= x"0000021a1";
		when x"00b11" => DOUT <= x"000002120";
		when x"00b12" => DOUT <= x"000202141";
		when x"00b13" => DOUT <= x"000202140";
		when x"00b14" => DOUT <= x"000003121";
		when x"00b15" => DOUT <= x"0000031a0";
		when x"00b16" => DOUT <= x"0002031c1";
		when x"00b17" => DOUT <= x"0002031c0";
		when x"00b18" => DOUT <= x"0000021a1";
		when x"00b19" => DOUT <= x"000002120";
		when x"00b1a" => DOUT <= x"000202141";
		when x"00b1b" => DOUT <= x"000202140";
		when x"00b1c" => DOUT <= x"000003121";
		when x"00b1d" => DOUT <= x"0000031a0";
		when x"00b1e" => DOUT <= x"0002031c1";
		when x"00b1f" => DOUT <= x"0002031c0";
		when x"00b20" => DOUT <= x"0000021a1";
		when x"00b21" => DOUT <= x"000002120";
		when x"00b22" => DOUT <= x"000202141";
		when x"00b23" => DOUT <= x"000202140";
		when x"00b24" => DOUT <= x"000003121";
		when x"00b25" => DOUT <= x"0000031a0";
		when x"00b26" => DOUT <= x"0002031c1";
		when x"00b27" => DOUT <= x"0002031c0";
		when x"00b28" => DOUT <= x"0000021a1";
		when x"00b29" => DOUT <= x"000002120";
		when x"00b2a" => DOUT <= x"000202141";
		when x"00b2b" => DOUT <= x"000202140";
		when x"00b2c" => DOUT <= x"000003121";
		when x"00b2d" => DOUT <= x"0000031a0";
		when x"00b2e" => DOUT <= x"0002031c1";
		when x"00b2f" => DOUT <= x"0002031c0";
		when x"00b30" => DOUT <= x"0000021a1";
		when x"00b31" => DOUT <= x"000002120";
		when x"00b32" => DOUT <= x"000202141";
		when x"00b33" => DOUT <= x"000202140";
		when x"00b34" => DOUT <= x"000003121";
		when x"00b35" => DOUT <= x"0000031a0";
		when x"00b36" => DOUT <= x"0002031c1";
		when x"00b37" => DOUT <= x"0002031c0";
		when x"00b38" => DOUT <= x"0000021a1";
		when x"00b39" => DOUT <= x"000002120";
		when x"00b3a" => DOUT <= x"000202141";
		when x"00b3b" => DOUT <= x"000202140";
		when x"00b3c" => DOUT <= x"000003121";
		when x"00b3d" => DOUT <= x"0000031a0";
		when x"00b3e" => DOUT <= x"0002031c1";
		when x"00b3f" => DOUT <= x"0002031c0";
		when x"00b40" => DOUT <= x"0000021a1";
		when x"00b41" => DOUT <= x"000002120";
		when x"00b42" => DOUT <= x"000202141";
		when x"00b43" => DOUT <= x"000202140";
		when x"00b44" => DOUT <= x"000003121";
		when x"00b45" => DOUT <= x"0000031a0";
		when x"00b46" => DOUT <= x"0002031c1";
		when x"00b47" => DOUT <= x"0002031c0";
		when x"00b48" => DOUT <= x"0000021a1";
		when x"00b49" => DOUT <= x"000002120";
		when x"00b4a" => DOUT <= x"000202141";
		when x"00b4b" => DOUT <= x"000202140";
		when x"00b4c" => DOUT <= x"000003121";
		when x"00b4d" => DOUT <= x"0000031a0";
		when x"00b4e" => DOUT <= x"0002031c1";
		when x"00b4f" => DOUT <= x"0002031c0";
		when x"00b50" => DOUT <= x"0000021a1";
		when x"00b51" => DOUT <= x"000002120";
		when x"00b52" => DOUT <= x"000202141";
		when x"00b53" => DOUT <= x"000202140";
		when x"00b54" => DOUT <= x"000003121";
		when x"00b55" => DOUT <= x"0000031a0";
		when x"00b56" => DOUT <= x"0002031c1";
		when x"00b57" => DOUT <= x"0002031c0";
		when x"00b58" => DOUT <= x"0000021a1";
		when x"00b59" => DOUT <= x"000002120";
		when x"00b5a" => DOUT <= x"000202141";
		when x"00b5b" => DOUT <= x"000202140";
		when x"00b5c" => DOUT <= x"000003121";
		when x"00b5d" => DOUT <= x"0000031a0";
		when x"00b5e" => DOUT <= x"0002031c1";
		when x"00b5f" => DOUT <= x"0002031c0";
		when x"00b60" => DOUT <= x"0000021a1";
		when x"00b61" => DOUT <= x"000002120";
		when x"00b62" => DOUT <= x"000202141";
		when x"00b63" => DOUT <= x"000202140";
		when x"00b64" => DOUT <= x"000003121";
		when x"00b65" => DOUT <= x"0000031a0";
		when x"00b66" => DOUT <= x"0002031c1";
		when x"00b67" => DOUT <= x"0002031c0";
		when x"00b68" => DOUT <= x"0000021a1";
		when x"00b69" => DOUT <= x"000002120";
		when x"00b6a" => DOUT <= x"000202141";
		when x"00b6b" => DOUT <= x"000202140";
		when x"00b6c" => DOUT <= x"000003121";
		when x"00b6d" => DOUT <= x"0000031a0";
		when x"00b6e" => DOUT <= x"0002031c1";
		when x"00b6f" => DOUT <= x"0002031c0";
		when x"00b70" => DOUT <= x"0000021a1";
		when x"00b71" => DOUT <= x"000002120";
		when x"00b72" => DOUT <= x"000202141";
		when x"00b73" => DOUT <= x"000202140";
		when x"00b74" => DOUT <= x"000003121";
		when x"00b75" => DOUT <= x"0000031a0";
		when x"00b76" => DOUT <= x"0002031c1";
		when x"00b77" => DOUT <= x"0002031c0";
		when x"00b78" => DOUT <= x"0000021a1";
		when x"00b79" => DOUT <= x"000002120";
		when x"00b7a" => DOUT <= x"000202141";
		when x"00b7b" => DOUT <= x"000202140";
		when x"00b7c" => DOUT <= x"000003121";
		when x"00b7d" => DOUT <= x"0000031a0";
		when x"00b7e" => DOUT <= x"0002031c1";
		when x"00b7f" => DOUT <= x"0002031c0";
		when x"00b80" => DOUT <= x"0000021a1";
		when x"00b81" => DOUT <= x"000002120";
		when x"00b82" => DOUT <= x"000202141";
		when x"00b83" => DOUT <= x"000202140";
		when x"00b84" => DOUT <= x"000003121";
		when x"00b85" => DOUT <= x"0000031a0";
		when x"00b86" => DOUT <= x"0002031c1";
		when x"00b87" => DOUT <= x"0002031c0";
		when x"00b88" => DOUT <= x"0000021a1";
		when x"00b89" => DOUT <= x"000002120";
		when x"00b8a" => DOUT <= x"000202141";
		when x"00b8b" => DOUT <= x"000202140";
		when x"00b8c" => DOUT <= x"000003121";
		when x"00b8d" => DOUT <= x"0000031a0";
		when x"00b8e" => DOUT <= x"0002031c1";
		when x"00b8f" => DOUT <= x"0002031c0";
		when x"00b90" => DOUT <= x"0000021a1";
		when x"00b91" => DOUT <= x"000002120";
		when x"00b92" => DOUT <= x"000202141";
		when x"00b93" => DOUT <= x"000202140";
		when x"00b94" => DOUT <= x"000003121";
		when x"00b95" => DOUT <= x"0000031a0";
		when x"00b96" => DOUT <= x"0002031c1";
		when x"00b97" => DOUT <= x"0002031c0";
		when x"00b98" => DOUT <= x"0000021a1";
		when x"00b99" => DOUT <= x"000002120";
		when x"00b9a" => DOUT <= x"000202141";
		when x"00b9b" => DOUT <= x"000202140";
		when x"00b9c" => DOUT <= x"000003121";
		when x"00b9d" => DOUT <= x"0000031a0";
		when x"00b9e" => DOUT <= x"0002031c1";
		when x"00b9f" => DOUT <= x"0002031c0";
		when x"00ba0" => DOUT <= x"0000021a1";
		when x"00ba1" => DOUT <= x"000002120";
		when x"00ba2" => DOUT <= x"000202141";
		when x"00ba3" => DOUT <= x"000202140";
		when x"00ba4" => DOUT <= x"000003121";
		when x"00ba5" => DOUT <= x"0000031a0";
		when x"00ba6" => DOUT <= x"0002031c1";
		when x"00ba7" => DOUT <= x"0002031c0";
		when x"00ba8" => DOUT <= x"0000021a1";
		when x"00ba9" => DOUT <= x"000002120";
		when x"00baa" => DOUT <= x"000202141";
		when x"00bab" => DOUT <= x"000202140";
		when x"00bac" => DOUT <= x"000003121";
		when x"00bad" => DOUT <= x"0000031a0";
		when x"00bae" => DOUT <= x"0002031c1";
		when x"00baf" => DOUT <= x"0002031c0";
		when x"00bb0" => DOUT <= x"0000021a1";
		when x"00bb1" => DOUT <= x"000002120";
		when x"00bb2" => DOUT <= x"000202141";
		when x"00bb3" => DOUT <= x"000202140";
		when x"00bb4" => DOUT <= x"000003121";
		when x"00bb5" => DOUT <= x"0000031a0";
		when x"00bb6" => DOUT <= x"0002031c1";
		when x"00bb7" => DOUT <= x"0002031c0";
		when x"00bb8" => DOUT <= x"0000021a1";
		when x"00bb9" => DOUT <= x"000002120";
		when x"00bba" => DOUT <= x"000202141";
		when x"00bbb" => DOUT <= x"000202140";
		when x"00bbc" => DOUT <= x"000003121";
		when x"00bbd" => DOUT <= x"0000031a0";
		when x"00bbe" => DOUT <= x"0002031c1";
		when x"00bbf" => DOUT <= x"0002031c0";
		when x"00bc0" => DOUT <= x"0000021a1";
		when x"00bc1" => DOUT <= x"000002120";
		when x"00bc2" => DOUT <= x"000202141";
		when x"00bc3" => DOUT <= x"000202140";
		when x"00bc4" => DOUT <= x"000003121";
		when x"00bc5" => DOUT <= x"0000031a0";
		when x"00bc6" => DOUT <= x"0002031c1";
		when x"00bc7" => DOUT <= x"0002031c0";
		when x"00bc8" => DOUT <= x"0000021a1";
		when x"00bc9" => DOUT <= x"000002120";
		when x"00bca" => DOUT <= x"000202141";
		when x"00bcb" => DOUT <= x"000202140";
		when x"00bcc" => DOUT <= x"000003121";
		when x"00bcd" => DOUT <= x"0000031a0";
		when x"00bce" => DOUT <= x"0002031c1";
		when x"00bcf" => DOUT <= x"0002031c0";
		when x"00bd0" => DOUT <= x"0000021a1";
		when x"00bd1" => DOUT <= x"000002120";
		when x"00bd2" => DOUT <= x"000202141";
		when x"00bd3" => DOUT <= x"000202140";
		when x"00bd4" => DOUT <= x"000003121";
		when x"00bd5" => DOUT <= x"0000031a0";
		when x"00bd6" => DOUT <= x"0002031c1";
		when x"00bd7" => DOUT <= x"0002031c0";
		when x"00bd8" => DOUT <= x"0000021a1";
		when x"00bd9" => DOUT <= x"000002120";
		when x"00bda" => DOUT <= x"000202141";
		when x"00bdb" => DOUT <= x"000202140";
		when x"00bdc" => DOUT <= x"000003121";
		when x"00bdd" => DOUT <= x"0000031a0";
		when x"00bde" => DOUT <= x"0002031c1";
		when x"00bdf" => DOUT <= x"0002031c0";
		when x"00be0" => DOUT <= x"0000021a1";
		when x"00be1" => DOUT <= x"000002120";
		when x"00be2" => DOUT <= x"000202141";
		when x"00be3" => DOUT <= x"000202140";
		when x"00be4" => DOUT <= x"000003121";
		when x"00be5" => DOUT <= x"0000031a0";
		when x"00be6" => DOUT <= x"0002031c1";
		when x"00be7" => DOUT <= x"0002031c0";
		when x"00be8" => DOUT <= x"0000021a1";
		when x"00be9" => DOUT <= x"000002120";
		when x"00bea" => DOUT <= x"000202141";
		when x"00beb" => DOUT <= x"000202140";
		when x"00bec" => DOUT <= x"000003121";
		when x"00bed" => DOUT <= x"0000031a0";
		when x"00bee" => DOUT <= x"0002031c1";
		when x"00bef" => DOUT <= x"0002031c0";
		when x"00bf0" => DOUT <= x"0000021a1";
		when x"00bf1" => DOUT <= x"000002120";
		when x"00bf2" => DOUT <= x"000202141";
		when x"00bf3" => DOUT <= x"000202140";
		when x"00bf4" => DOUT <= x"000003121";
		when x"00bf5" => DOUT <= x"0000031a0";
		when x"00bf6" => DOUT <= x"0002031c1";
		when x"00bf7" => DOUT <= x"0002031c0";
		when x"00bf8" => DOUT <= x"0000021a1";
		when x"00bf9" => DOUT <= x"000002120";
		when x"00bfa" => DOUT <= x"000202141";
		when x"00bfb" => DOUT <= x"000202140";
		when x"00bfc" => DOUT <= x"000003121";
		when x"00bfd" => DOUT <= x"0000031a0";
		when x"00bfe" => DOUT <= x"0002031c1";
		when x"00bff" => DOUT <= x"0002031c0";
		when x"00c00" => DOUT <= x"0000021a1";
		when x"00c01" => DOUT <= x"000002120";
		when x"00c02" => DOUT <= x"000202141";
		when x"00c03" => DOUT <= x"000202140";
		when x"00c04" => DOUT <= x"000003121";
		when x"00c05" => DOUT <= x"0000031a0";
		when x"00c06" => DOUT <= x"0002031c1";
		when x"00c07" => DOUT <= x"0002031c0";
		when x"00c08" => DOUT <= x"0000021a1";
		when x"00c09" => DOUT <= x"000002120";
		when x"00c0a" => DOUT <= x"000202141";
		when x"00c0b" => DOUT <= x"000202140";
		when x"00c0c" => DOUT <= x"000003121";
		when x"00c0d" => DOUT <= x"0000031a0";
		when x"00c0e" => DOUT <= x"0002031c1";
		when x"00c0f" => DOUT <= x"0002031c0";
		when x"00c10" => DOUT <= x"0000021a1";
		when x"00c11" => DOUT <= x"000002120";
		when x"00c12" => DOUT <= x"000202141";
		when x"00c13" => DOUT <= x"000202140";
		when x"00c14" => DOUT <= x"000003121";
		when x"00c15" => DOUT <= x"0000031a0";
		when x"00c16" => DOUT <= x"0002031c1";
		when x"00c17" => DOUT <= x"0002031c0";
		when x"00c18" => DOUT <= x"0000021a1";
		when x"00c19" => DOUT <= x"000002120";
		when x"00c1a" => DOUT <= x"000202141";
		when x"00c1b" => DOUT <= x"000202140";
		when x"00c1c" => DOUT <= x"000003121";
		when x"00c1d" => DOUT <= x"0000031a0";
		when x"00c1e" => DOUT <= x"0002031c1";
		when x"00c1f" => DOUT <= x"0002031c0";
		when x"00c20" => DOUT <= x"0000021a1";
		when x"00c21" => DOUT <= x"000002120";
		when x"00c22" => DOUT <= x"000202141";
		when x"00c23" => DOUT <= x"000202140";
		when x"00c24" => DOUT <= x"000003121";
		when x"00c25" => DOUT <= x"0000031a0";
		when x"00c26" => DOUT <= x"0002031c1";
		when x"00c27" => DOUT <= x"0002031c0";
		when x"00c28" => DOUT <= x"0000021a1";
		when x"00c29" => DOUT <= x"000002120";
		when x"00c2a" => DOUT <= x"000202141";
		when x"00c2b" => DOUT <= x"000202140";
		when x"00c2c" => DOUT <= x"000003121";
		when x"00c2d" => DOUT <= x"0000031a0";
		when x"00c2e" => DOUT <= x"0002031c1";
		when x"00c2f" => DOUT <= x"0002031c0";
		when x"00c30" => DOUT <= x"0000021a1";
		when x"00c31" => DOUT <= x"000002120";
		when x"00c32" => DOUT <= x"000202141";
		when x"00c33" => DOUT <= x"000202140";
		when x"00c34" => DOUT <= x"000003121";
		when x"00c35" => DOUT <= x"0000031a0";
		when x"00c36" => DOUT <= x"0002031c1";
		when x"00c37" => DOUT <= x"0002031c0";
		when x"00c38" => DOUT <= x"0000021a1";
		when x"00c39" => DOUT <= x"000002120";
		when x"00c3a" => DOUT <= x"000202141";
		when x"00c3b" => DOUT <= x"000202140";
		when x"00c3c" => DOUT <= x"000003121";
		when x"00c3d" => DOUT <= x"0000031a0";
		when x"00c3e" => DOUT <= x"0002031c1";
		when x"00c3f" => DOUT <= x"0002031c0";
		when x"00c40" => DOUT <= x"0000021a1";
		when x"00c41" => DOUT <= x"000002120";
		when x"00c42" => DOUT <= x"000202141";
		when x"00c43" => DOUT <= x"000202140";
		when x"00c44" => DOUT <= x"000003121";
		when x"00c45" => DOUT <= x"0000031a0";
		when x"00c46" => DOUT <= x"0002031c1";
		when x"00c47" => DOUT <= x"0002031c0";
		when x"00c48" => DOUT <= x"0000021a1";
		when x"00c49" => DOUT <= x"000002120";
		when x"00c4a" => DOUT <= x"000202141";
		when x"00c4b" => DOUT <= x"000202140";
		when x"00c4c" => DOUT <= x"000003121";
		when x"00c4d" => DOUT <= x"0000031a0";
		when x"00c4e" => DOUT <= x"0002031c1";
		when x"00c4f" => DOUT <= x"0002031c0";
		when x"00c50" => DOUT <= x"0000021a1";
		when x"00c51" => DOUT <= x"000002120";
		when x"00c52" => DOUT <= x"000202141";
		when x"00c53" => DOUT <= x"000202140";
		when x"00c54" => DOUT <= x"000003121";
		when x"00c55" => DOUT <= x"0000031a0";
		when x"00c56" => DOUT <= x"0002031c1";
		when x"00c57" => DOUT <= x"0002031c0";
		when x"00c58" => DOUT <= x"0000021a1";
		when x"00c59" => DOUT <= x"000002120";
		when x"00c5a" => DOUT <= x"000202141";
		when x"00c5b" => DOUT <= x"000202140";
		when x"00c5c" => DOUT <= x"000003121";
		when x"00c5d" => DOUT <= x"0000031a0";
		when x"00c5e" => DOUT <= x"0002031c1";
		when x"00c5f" => DOUT <= x"0002031c0";
		when x"00c60" => DOUT <= x"0000021a1";
		when x"00c61" => DOUT <= x"000002120";
		when x"00c62" => DOUT <= x"000202141";
		when x"00c63" => DOUT <= x"000202140";
		when x"00c64" => DOUT <= x"000003121";
		when x"00c65" => DOUT <= x"0000031a0";
		when x"00c66" => DOUT <= x"0002031c1";
		when x"00c67" => DOUT <= x"0002031c0";
		when x"00c68" => DOUT <= x"0000021a1";
		when x"00c69" => DOUT <= x"000002120";
		when x"00c6a" => DOUT <= x"000202141";
		when x"00c6b" => DOUT <= x"000202140";
		when x"00c6c" => DOUT <= x"000003121";
		when x"00c6d" => DOUT <= x"0000031a0";
		when x"00c6e" => DOUT <= x"0002031c1";
		when x"00c6f" => DOUT <= x"0002031c0";
		when x"00c70" => DOUT <= x"0000021a1";
		when x"00c71" => DOUT <= x"000002120";
		when x"00c72" => DOUT <= x"000202141";
		when x"00c73" => DOUT <= x"000202140";
		when x"00c74" => DOUT <= x"000003121";
		when x"00c75" => DOUT <= x"0000031a0";
		when x"00c76" => DOUT <= x"0002031c1";
		when x"00c77" => DOUT <= x"0002031c0";
		when x"00c78" => DOUT <= x"0000021a1";
		when x"00c79" => DOUT <= x"000002120";
		when x"00c7a" => DOUT <= x"000202141";
		when x"00c7b" => DOUT <= x"000202140";
		when x"00c7c" => DOUT <= x"000003121";
		when x"00c7d" => DOUT <= x"0000031a0";
		when x"00c7e" => DOUT <= x"0002031c1";
		when x"00c7f" => DOUT <= x"0002031c0";
		when x"00c80" => DOUT <= x"0000021a1";
		when x"00c81" => DOUT <= x"000002120";
		when x"00c82" => DOUT <= x"000202141";
		when x"00c83" => DOUT <= x"000202140";
		when x"00c84" => DOUT <= x"000003121";
		when x"00c85" => DOUT <= x"0000031a0";
		when x"00c86" => DOUT <= x"0002031c1";
		when x"00c87" => DOUT <= x"0002031c0";
		when x"00c88" => DOUT <= x"0000021a1";
		when x"00c89" => DOUT <= x"000002120";
		when x"00c8a" => DOUT <= x"000202141";
		when x"00c8b" => DOUT <= x"000202140";
		when x"00c8c" => DOUT <= x"000003121";
		when x"00c8d" => DOUT <= x"0000031a0";
		when x"00c8e" => DOUT <= x"0002031c1";
		when x"00c8f" => DOUT <= x"0002031c0";
		when x"00c90" => DOUT <= x"0000021a1";
		when x"00c91" => DOUT <= x"000002120";
		when x"00c92" => DOUT <= x"000202141";
		when x"00c93" => DOUT <= x"000202140";
		when x"00c94" => DOUT <= x"000003121";
		when x"00c95" => DOUT <= x"0000031a0";
		when x"00c96" => DOUT <= x"0002031c1";
		when x"00c97" => DOUT <= x"0002031c0";
		when x"00c98" => DOUT <= x"0000021a1";
		when x"00c99" => DOUT <= x"000002120";
		when x"00c9a" => DOUT <= x"000202141";
		when x"00c9b" => DOUT <= x"000202140";
		when x"00c9c" => DOUT <= x"000003121";
		when x"00c9d" => DOUT <= x"0000031a0";
		when x"00c9e" => DOUT <= x"0002031c1";
		when x"00c9f" => DOUT <= x"0002031c0";
		when x"00ca0" => DOUT <= x"0000021a1";
		when x"00ca1" => DOUT <= x"000002120";
		when x"00ca2" => DOUT <= x"000202141";
		when x"00ca3" => DOUT <= x"000202140";
		when x"00ca4" => DOUT <= x"000003121";
		when x"00ca5" => DOUT <= x"0000031a0";
		when x"00ca6" => DOUT <= x"0002031c1";
		when x"00ca7" => DOUT <= x"0002031c0";
		when x"00ca8" => DOUT <= x"0000021a1";
		when x"00ca9" => DOUT <= x"000002120";
		when x"00caa" => DOUT <= x"000202141";
		when x"00cab" => DOUT <= x"000202140";
		when x"00cac" => DOUT <= x"000003121";
		when x"00cad" => DOUT <= x"0000031a0";
		when x"00cae" => DOUT <= x"0002031c1";
		when x"00caf" => DOUT <= x"0002031c0";
		when x"00cb0" => DOUT <= x"0000021a1";
		when x"00cb1" => DOUT <= x"000002120";
		when x"00cb2" => DOUT <= x"000202141";
		when x"00cb3" => DOUT <= x"000202140";
		when x"00cb4" => DOUT <= x"000003121";
		when x"00cb5" => DOUT <= x"0000031a0";
		when x"00cb6" => DOUT <= x"0002031c1";
		when x"00cb7" => DOUT <= x"0002031c0";
		when x"00cb8" => DOUT <= x"0000021a1";
		when x"00cb9" => DOUT <= x"000002120";
		when x"00cba" => DOUT <= x"000202141";
		when x"00cbb" => DOUT <= x"000202140";
		when x"00cbc" => DOUT <= x"000003121";
		when x"00cbd" => DOUT <= x"0000031a0";
		when x"00cbe" => DOUT <= x"0002031c1";
		when x"00cbf" => DOUT <= x"0002031c0";
		when x"00cc0" => DOUT <= x"0000021a1";
		when x"00cc1" => DOUT <= x"000002120";
		when x"00cc2" => DOUT <= x"000202141";
		when x"00cc3" => DOUT <= x"000202140";
		when x"00cc4" => DOUT <= x"000003121";
		when x"00cc5" => DOUT <= x"0000031a0";
		when x"00cc6" => DOUT <= x"0002031c1";
		when x"00cc7" => DOUT <= x"0002031c0";
		when x"00cc8" => DOUT <= x"0000021a1";
		when x"00cc9" => DOUT <= x"000002120";
		when x"00cca" => DOUT <= x"000202141";
		when x"00ccb" => DOUT <= x"000202140";
		when x"00ccc" => DOUT <= x"000003121";
		when x"00ccd" => DOUT <= x"0000031a0";
		when x"00cce" => DOUT <= x"0002031c1";
		when x"00ccf" => DOUT <= x"0002031c0";
		when x"00cd0" => DOUT <= x"0000021a1";
		when x"00cd1" => DOUT <= x"000002120";
		when x"00cd2" => DOUT <= x"000202141";
		when x"00cd3" => DOUT <= x"000202140";
		when x"00cd4" => DOUT <= x"000003121";
		when x"00cd5" => DOUT <= x"0000031a0";
		when x"00cd6" => DOUT <= x"0002031c1";
		when x"00cd7" => DOUT <= x"0002031c0";
		when x"00cd8" => DOUT <= x"0000021a1";
		when x"00cd9" => DOUT <= x"000002120";
		when x"00cda" => DOUT <= x"000202141";
		when x"00cdb" => DOUT <= x"000202140";
		when x"00cdc" => DOUT <= x"000003121";
		when x"00cdd" => DOUT <= x"0000031a0";
		when x"00cde" => DOUT <= x"0002031c1";
		when x"00cdf" => DOUT <= x"0002031c0";
		when x"00ce0" => DOUT <= x"0000021a1";
		when x"00ce1" => DOUT <= x"000002120";
		when x"00ce2" => DOUT <= x"000202141";
		when x"00ce3" => DOUT <= x"000202140";
		when x"00ce4" => DOUT <= x"000003121";
		when x"00ce5" => DOUT <= x"0000031a0";
		when x"00ce6" => DOUT <= x"0002031c1";
		when x"00ce7" => DOUT <= x"0002031c0";
		when x"00ce8" => DOUT <= x"0000021a1";
		when x"00ce9" => DOUT <= x"000002120";
		when x"00cea" => DOUT <= x"000202141";
		when x"00ceb" => DOUT <= x"000202140";
		when x"00cec" => DOUT <= x"000003121";
		when x"00ced" => DOUT <= x"0000031a0";
		when x"00cee" => DOUT <= x"0002031c1";
		when x"00cef" => DOUT <= x"0002031c0";
		when x"00cf0" => DOUT <= x"0000021a1";
		when x"00cf1" => DOUT <= x"000002120";
		when x"00cf2" => DOUT <= x"000202141";
		when x"00cf3" => DOUT <= x"000202140";
		when x"00cf4" => DOUT <= x"000003121";
		when x"00cf5" => DOUT <= x"0000031a0";
		when x"00cf6" => DOUT <= x"0002031c1";
		when x"00cf7" => DOUT <= x"0002031c0";
		when x"00cf8" => DOUT <= x"0000021a1";
		when x"00cf9" => DOUT <= x"000002120";
		when x"00cfa" => DOUT <= x"000202141";
		when x"00cfb" => DOUT <= x"000202140";
		when x"00cfc" => DOUT <= x"000003121";
		when x"00cfd" => DOUT <= x"0000031a0";
		when x"00cfe" => DOUT <= x"0002031c1";
		when x"00cff" => DOUT <= x"0002031c0";
		when x"00d00" => DOUT <= x"0000021a1";
		when x"00d01" => DOUT <= x"000002120";
		when x"00d02" => DOUT <= x"000202141";
		when x"00d03" => DOUT <= x"000202140";
		when x"00d04" => DOUT <= x"000003121";
		when x"00d05" => DOUT <= x"0000031a0";
		when x"00d06" => DOUT <= x"0002031c1";
		when x"00d07" => DOUT <= x"0002031c0";
		when x"00d08" => DOUT <= x"0000021a1";
		when x"00d09" => DOUT <= x"000002120";
		when x"00d0a" => DOUT <= x"000202141";
		when x"00d0b" => DOUT <= x"000202140";
		when x"00d0c" => DOUT <= x"000003121";
		when x"00d0d" => DOUT <= x"0000031a0";
		when x"00d0e" => DOUT <= x"0002031c1";
		when x"00d0f" => DOUT <= x"0002031c0";
		when x"00d10" => DOUT <= x"0000021a1";
		when x"00d11" => DOUT <= x"000002120";
		when x"00d12" => DOUT <= x"000202141";
		when x"00d13" => DOUT <= x"000202140";
		when x"00d14" => DOUT <= x"000003121";
		when x"00d15" => DOUT <= x"0000031a0";
		when x"00d16" => DOUT <= x"0002031c1";
		when x"00d17" => DOUT <= x"0002031c0";
		when x"00d18" => DOUT <= x"0000021a1";
		when x"00d19" => DOUT <= x"000002120";
		when x"00d1a" => DOUT <= x"000202141";
		when x"00d1b" => DOUT <= x"000202140";
		when x"00d1c" => DOUT <= x"000003121";
		when x"00d1d" => DOUT <= x"0000031a0";
		when x"00d1e" => DOUT <= x"0002031c1";
		when x"00d1f" => DOUT <= x"0002031c0";
		when x"00d20" => DOUT <= x"0000021a1";
		when x"00d21" => DOUT <= x"000002120";
		when x"00d22" => DOUT <= x"000202141";
		when x"00d23" => DOUT <= x"000202140";
		when x"00d24" => DOUT <= x"000003121";
		when x"00d25" => DOUT <= x"0000031a0";
		when x"00d26" => DOUT <= x"0002031c1";
		when x"00d27" => DOUT <= x"0002031c0";
		when x"00d28" => DOUT <= x"0000021a1";
		when x"00d29" => DOUT <= x"000002120";
		when x"00d2a" => DOUT <= x"000202141";
		when x"00d2b" => DOUT <= x"000202140";
		when x"00d2c" => DOUT <= x"000003121";
		when x"00d2d" => DOUT <= x"0000031a0";
		when x"00d2e" => DOUT <= x"0002031c1";
		when x"00d2f" => DOUT <= x"0002031c0";
		when x"00d30" => DOUT <= x"0000021a1";
		when x"00d31" => DOUT <= x"000002120";
		when x"00d32" => DOUT <= x"000202141";
		when x"00d33" => DOUT <= x"000202140";
		when x"00d34" => DOUT <= x"000003121";
		when x"00d35" => DOUT <= x"0000031a0";
		when x"00d36" => DOUT <= x"0002031c1";
		when x"00d37" => DOUT <= x"0002031c0";
		when x"00d38" => DOUT <= x"0000021a1";
		when x"00d39" => DOUT <= x"000002120";
		when x"00d3a" => DOUT <= x"000202141";
		when x"00d3b" => DOUT <= x"000202140";
		when x"00d3c" => DOUT <= x"000003121";
		when x"00d3d" => DOUT <= x"0000031a0";
		when x"00d3e" => DOUT <= x"0002031c1";
		when x"00d3f" => DOUT <= x"0002031c0";
		when x"00d40" => DOUT <= x"0000021a1";
		when x"00d41" => DOUT <= x"000002120";
		when x"00d42" => DOUT <= x"000202141";
		when x"00d43" => DOUT <= x"000202140";
		when x"00d44" => DOUT <= x"000003121";
		when x"00d45" => DOUT <= x"0000031a0";
		when x"00d46" => DOUT <= x"0002031c1";
		when x"00d47" => DOUT <= x"0002031c0";
		when x"00d48" => DOUT <= x"0000021a1";
		when x"00d49" => DOUT <= x"000002120";
		when x"00d4a" => DOUT <= x"000202141";
		when x"00d4b" => DOUT <= x"000202140";
		when x"00d4c" => DOUT <= x"000003121";
		when x"00d4d" => DOUT <= x"0000031a0";
		when x"00d4e" => DOUT <= x"0002031c1";
		when x"00d4f" => DOUT <= x"0002031c0";
		when x"00d50" => DOUT <= x"0000021a1";
		when x"00d51" => DOUT <= x"000002120";
		when x"00d52" => DOUT <= x"000202141";
		when x"00d53" => DOUT <= x"000202140";
		when x"00d54" => DOUT <= x"000003121";
		when x"00d55" => DOUT <= x"0000031a0";
		when x"00d56" => DOUT <= x"0002031c1";
		when x"00d57" => DOUT <= x"0002031c0";
		when x"00d58" => DOUT <= x"0000021a1";
		when x"00d59" => DOUT <= x"000002120";
		when x"00d5a" => DOUT <= x"000202141";
		when x"00d5b" => DOUT <= x"000202140";
		when x"00d5c" => DOUT <= x"000003121";
		when x"00d5d" => DOUT <= x"0000031a0";
		when x"00d5e" => DOUT <= x"0002031c1";
		when x"00d5f" => DOUT <= x"0002031c0";
		when x"00d60" => DOUT <= x"0000021a1";
		when x"00d61" => DOUT <= x"000002120";
		when x"00d62" => DOUT <= x"000202141";
		when x"00d63" => DOUT <= x"000202140";
		when x"00d64" => DOUT <= x"000003121";
		when x"00d65" => DOUT <= x"0000031a0";
		when x"00d66" => DOUT <= x"0002031c1";
		when x"00d67" => DOUT <= x"0002031c0";
		when x"00d68" => DOUT <= x"0000021a1";
		when x"00d69" => DOUT <= x"000002120";
		when x"00d6a" => DOUT <= x"000202141";
		when x"00d6b" => DOUT <= x"000202140";
		when x"00d6c" => DOUT <= x"000003121";
		when x"00d6d" => DOUT <= x"0000031a0";
		when x"00d6e" => DOUT <= x"0002031c1";
		when x"00d6f" => DOUT <= x"0002031c0";
		when x"00d70" => DOUT <= x"0000001a1";
		when x"00d71" => DOUT <= x"000000120";
		when x"00d72" => DOUT <= x"000200141";
		when x"00d73" => DOUT <= x"000200140";
		when x"00d74" => DOUT <= x"000001121";
		when x"00d75" => DOUT <= x"0000011a0";
		when x"00d76" => DOUT <= x"0002011c1";
		when x"00d77" => DOUT <= x"0002011c0";
		when x"00d78" => DOUT <= x"0000001a1";
		when x"00d79" => DOUT <= x"000000120";
		when x"00d7a" => DOUT <= x"000200141";
		when x"00d7b" => DOUT <= x"000200140";
		when x"00d7c" => DOUT <= x"000001121";
		when x"00d7d" => DOUT <= x"0000011a0";
		when x"00d7e" => DOUT <= x"0002011c1";
		when x"00d7f" => DOUT <= x"0002011c0";
		when x"00d80" => DOUT <= x"0000021a1";
		when x"00d81" => DOUT <= x"000002120";
		when x"00d82" => DOUT <= x"000202141";
		when x"00d83" => DOUT <= x"000202140";
		when x"00d84" => DOUT <= x"000003121";
		when x"00d85" => DOUT <= x"0000031a0";
		when x"00d86" => DOUT <= x"0002031c1";
		when x"00d87" => DOUT <= x"0002031c0";
		when x"00d88" => DOUT <= x"0000021a1";
		when x"00d89" => DOUT <= x"000002120";
		when x"00d8a" => DOUT <= x"000202141";
		when x"00d8b" => DOUT <= x"000202140";
		when x"00d8c" => DOUT <= x"000003121";
		when x"00d8d" => DOUT <= x"0000031a0";
		when x"00d8e" => DOUT <= x"0002031c1";
		when x"00d8f" => DOUT <= x"0002031c0";
		when x"00d90" => DOUT <= x"0000021a1";
		when x"00d91" => DOUT <= x"000002120";
		when x"00d92" => DOUT <= x"000202141";
		when x"00d93" => DOUT <= x"000202140";
		when x"00d94" => DOUT <= x"000003121";
		when x"00d95" => DOUT <= x"0000031a0";
		when x"00d96" => DOUT <= x"0002031c1";
		when x"00d97" => DOUT <= x"0002031c0";
		when x"00d98" => DOUT <= x"0000021a1";
		when x"00d99" => DOUT <= x"000002120";
		when x"00d9a" => DOUT <= x"000202141";
		when x"00d9b" => DOUT <= x"000202140";
		when x"00d9c" => DOUT <= x"000003121";
		when x"00d9d" => DOUT <= x"0000031a0";
		when x"00d9e" => DOUT <= x"0002031c1";
		when x"00d9f" => DOUT <= x"0002031c0";
		when x"00da0" => DOUT <= x"0000021a1";
		when x"00da1" => DOUT <= x"000002120";
		when x"00da2" => DOUT <= x"000202141";
		when x"00da3" => DOUT <= x"000202140";
		when x"00da4" => DOUT <= x"000003121";
		when x"00da5" => DOUT <= x"0000031a0";
		when x"00da6" => DOUT <= x"0002031c1";
		when x"00da7" => DOUT <= x"0002031c0";
		when x"00da8" => DOUT <= x"0000021a1";
		when x"00da9" => DOUT <= x"000002120";
		when x"00daa" => DOUT <= x"000202141";
		when x"00dab" => DOUT <= x"000202140";
		when x"00dac" => DOUT <= x"000003121";
		when x"00dad" => DOUT <= x"0000031a0";
		when x"00dae" => DOUT <= x"0002031c1";
		when x"00daf" => DOUT <= x"0002031c0";
		when x"00db0" => DOUT <= x"0000001a1";
		when x"00db1" => DOUT <= x"000000120";
		when x"00db2" => DOUT <= x"000200141";
		when x"00db3" => DOUT <= x"000200140";
		when x"00db4" => DOUT <= x"000001121";
		when x"00db5" => DOUT <= x"0000011a0";
		when x"00db6" => DOUT <= x"0002011c1";
		when x"00db7" => DOUT <= x"0002011c0";
		when x"00db8" => DOUT <= x"0000001a1";
		when x"00db9" => DOUT <= x"000000120";
		when x"00dba" => DOUT <= x"000200141";
		when x"00dbb" => DOUT <= x"000200140";
		when x"00dbc" => DOUT <= x"000001121";
		when x"00dbd" => DOUT <= x"0000011a0";
		when x"00dbe" => DOUT <= x"0002011c1";
		when x"00dbf" => DOUT <= x"0002011c0";
		when x"00dc0" => DOUT <= x"0000021a1";
		when x"00dc1" => DOUT <= x"000002120";
		when x"00dc2" => DOUT <= x"000202141";
		when x"00dc3" => DOUT <= x"000202140";
		when x"00dc4" => DOUT <= x"000002121";
		when x"00dc5" => DOUT <= x"0000021a0";
		when x"00dc6" => DOUT <= x"0002021c1";
		when x"00dc7" => DOUT <= x"0002021c0";
		when x"00dc8" => DOUT <= x"0000021a1";
		when x"00dc9" => DOUT <= x"000002120";
		when x"00dca" => DOUT <= x"000202141";
		when x"00dcb" => DOUT <= x"000202140";
		when x"00dcc" => DOUT <= x"000002121";
		when x"00dcd" => DOUT <= x"0000021a0";
		when x"00dce" => DOUT <= x"0002021c1";
		when x"00dcf" => DOUT <= x"0002021c0";
		when x"00dd0" => DOUT <= x"0000021a1";
		when x"00dd1" => DOUT <= x"000002120";
		when x"00dd2" => DOUT <= x"000202141";
		when x"00dd3" => DOUT <= x"000202140";
		when x"00dd4" => DOUT <= x"000002121";
		when x"00dd5" => DOUT <= x"0000021a0";
		when x"00dd6" => DOUT <= x"0002021c1";
		when x"00dd7" => DOUT <= x"0002021c0";
		when x"00dd8" => DOUT <= x"0000021a1";
		when x"00dd9" => DOUT <= x"000002120";
		when x"00dda" => DOUT <= x"000202141";
		when x"00ddb" => DOUT <= x"000202140";
		when x"00ddc" => DOUT <= x"000002121";
		when x"00ddd" => DOUT <= x"0000021a0";
		when x"00dde" => DOUT <= x"0002021c1";
		when x"00ddf" => DOUT <= x"0002021c0";
		when x"00de0" => DOUT <= x"00001a1a1";
		when x"00de1" => DOUT <= x"00001a120";
		when x"00de2" => DOUT <= x"00021a141";
		when x"00de3" => DOUT <= x"00021a140";
		when x"00de4" => DOUT <= x"00001a121";
		when x"00de5" => DOUT <= x"00001a1a0";
		when x"00de6" => DOUT <= x"00021a1c1";
		when x"00de7" => DOUT <= x"00021a1c0";
		when x"00de8" => DOUT <= x"00001a1a1";
		when x"00de9" => DOUT <= x"00001a120";
		when x"00dea" => DOUT <= x"00021a141";
		when x"00deb" => DOUT <= x"00021a140";
		when x"00dec" => DOUT <= x"00001a121";
		when x"00ded" => DOUT <= x"00001a1a0";
		when x"00dee" => DOUT <= x"00021a1c1";
		when x"00def" => DOUT <= x"00021a1c0";
		when x"00df0" => DOUT <= x"00001a1a1";
		when x"00df1" => DOUT <= x"00001a120";
		when x"00df2" => DOUT <= x"00021a141";
		when x"00df3" => DOUT <= x"00021a140";
		when x"00df4" => DOUT <= x"00001a121";
		when x"00df5" => DOUT <= x"00001a1a0";
		when x"00df6" => DOUT <= x"00021a1c1";
		when x"00df7" => DOUT <= x"00021a1c0";
		when x"00df8" => DOUT <= x"00001a1a1";
		when x"00df9" => DOUT <= x"00001a120";
		when x"00dfa" => DOUT <= x"00021a141";
		when x"00dfb" => DOUT <= x"00021a140";
		when x"00dfc" => DOUT <= x"00001a121";
		when x"00dfd" => DOUT <= x"00001a1a0";
		when x"00dfe" => DOUT <= x"00021a1c1";
		when x"00dff" => DOUT <= x"00021a1c0";
		when x"00e00" => DOUT <= x"0000021a1";
		when x"00e01" => DOUT <= x"000002120";
		when x"00e02" => DOUT <= x"000202141";
		when x"00e03" => DOUT <= x"000202140";
		when x"00e04" => DOUT <= x"000002121";
		when x"00e05" => DOUT <= x"0000021a0";
		when x"00e06" => DOUT <= x"0002021c1";
		when x"00e07" => DOUT <= x"0002021c0";
		when x"00e08" => DOUT <= x"0000021a1";
		when x"00e09" => DOUT <= x"000002120";
		when x"00e0a" => DOUT <= x"000202141";
		when x"00e0b" => DOUT <= x"000202140";
		when x"00e0c" => DOUT <= x"000002121";
		when x"00e0d" => DOUT <= x"0000021a0";
		when x"00e0e" => DOUT <= x"0002021c1";
		when x"00e0f" => DOUT <= x"0002021c0";
		when x"00e10" => DOUT <= x"0000021a1";
		when x"00e11" => DOUT <= x"000002120";
		when x"00e12" => DOUT <= x"000202141";
		when x"00e13" => DOUT <= x"000202140";
		when x"00e14" => DOUT <= x"000002121";
		when x"00e15" => DOUT <= x"0000021a0";
		when x"00e16" => DOUT <= x"0002021c1";
		when x"00e17" => DOUT <= x"0002021c0";
		when x"00e18" => DOUT <= x"0000021a1";
		when x"00e19" => DOUT <= x"000002120";
		when x"00e1a" => DOUT <= x"000202141";
		when x"00e1b" => DOUT <= x"000202140";
		when x"00e1c" => DOUT <= x"000002121";
		when x"00e1d" => DOUT <= x"0000021a0";
		when x"00e1e" => DOUT <= x"0002021c1";
		when x"00e1f" => DOUT <= x"0002021c0";
		when x"00e20" => DOUT <= x"0000021a1";
		when x"00e21" => DOUT <= x"000002120";
		when x"00e22" => DOUT <= x"000202141";
		when x"00e23" => DOUT <= x"000202140";
		when x"00e24" => DOUT <= x"000002121";
		when x"00e25" => DOUT <= x"0000021a0";
		when x"00e26" => DOUT <= x"0002021c1";
		when x"00e27" => DOUT <= x"0002021c0";
		when x"00e28" => DOUT <= x"0000021a1";
		when x"00e29" => DOUT <= x"000002120";
		when x"00e2a" => DOUT <= x"000202141";
		when x"00e2b" => DOUT <= x"000202140";
		when x"00e2c" => DOUT <= x"000002121";
		when x"00e2d" => DOUT <= x"0000021a0";
		when x"00e2e" => DOUT <= x"0002021c1";
		when x"00e2f" => DOUT <= x"0002021c0";
		when x"00e30" => DOUT <= x"0000120a1";
		when x"00e31" => DOUT <= x"000012020";
		when x"00e32" => DOUT <= x"000212041";
		when x"00e33" => DOUT <= x"000212040";
		when x"00e34" => DOUT <= x"000012021";
		when x"00e35" => DOUT <= x"0000120a0";
		when x"00e36" => DOUT <= x"0002120c1";
		when x"00e37" => DOUT <= x"0002120c0";
		when x"00e38" => DOUT <= x"0000120a1";
		when x"00e39" => DOUT <= x"000012020";
		when x"00e3a" => DOUT <= x"000212041";
		when x"00e3b" => DOUT <= x"000212040";
		when x"00e3c" => DOUT <= x"000012021";
		when x"00e3d" => DOUT <= x"0000120a0";
		when x"00e3e" => DOUT <= x"0002120c1";
		when x"00e3f" => DOUT <= x"0002120c0";
		when x"00e40" => DOUT <= x"0000120a1";
		when x"00e41" => DOUT <= x"000012020";
		when x"00e42" => DOUT <= x"000212041";
		when x"00e43" => DOUT <= x"000212040";
		when x"00e44" => DOUT <= x"000012021";
		when x"00e45" => DOUT <= x"0000120a0";
		when x"00e46" => DOUT <= x"0002120c1";
		when x"00e47" => DOUT <= x"0002120c0";
		when x"00e48" => DOUT <= x"0000120a1";
		when x"00e49" => DOUT <= x"000012020";
		when x"00e4a" => DOUT <= x"000212041";
		when x"00e4b" => DOUT <= x"000212040";
		when x"00e4c" => DOUT <= x"000012021";
		when x"00e4d" => DOUT <= x"0000120a0";
		when x"00e4e" => DOUT <= x"0002120c1";
		when x"00e4f" => DOUT <= x"0002120c0";
		when x"00e50" => DOUT <= x"0000024a1";
		when x"00e51" => DOUT <= x"000002420";
		when x"00e52" => DOUT <= x"000202441";
		when x"00e53" => DOUT <= x"000202440";
		when x"00e54" => DOUT <= x"000002421";
		when x"00e55" => DOUT <= x"0000024a0";
		when x"00e56" => DOUT <= x"0002024c1";
		when x"00e57" => DOUT <= x"0002024c0";
		when x"00e58" => DOUT <= x"0000024a1";
		when x"00e59" => DOUT <= x"000002420";
		when x"00e5a" => DOUT <= x"000202441";
		when x"00e5b" => DOUT <= x"000202440";
		when x"00e5c" => DOUT <= x"000002421";
		when x"00e5d" => DOUT <= x"0000024a0";
		when x"00e5e" => DOUT <= x"0002024c1";
		when x"00e5f" => DOUT <= x"0002024c0";
		when x"00e60" => DOUT <= x"0000024a1";
		when x"00e61" => DOUT <= x"000002420";
		when x"00e62" => DOUT <= x"000202441";
		when x"00e63" => DOUT <= x"000202440";
		when x"00e64" => DOUT <= x"000002421";
		when x"00e65" => DOUT <= x"0000024a0";
		when x"00e66" => DOUT <= x"0002024c1";
		when x"00e67" => DOUT <= x"0002024c0";
		when x"00e68" => DOUT <= x"0000024a1";
		when x"00e69" => DOUT <= x"000002420";
		when x"00e6a" => DOUT <= x"000202441";
		when x"00e6b" => DOUT <= x"000202440";
		when x"00e6c" => DOUT <= x"000002421";
		when x"00e6d" => DOUT <= x"0000024a0";
		when x"00e6e" => DOUT <= x"0002024c1";
		when x"00e6f" => DOUT <= x"0002024c0";
		when x"00e70" => DOUT <= x"0000125a1";
		when x"00e71" => DOUT <= x"000012520";
		when x"00e72" => DOUT <= x"000212541";
		when x"00e73" => DOUT <= x"000212540";
		when x"00e74" => DOUT <= x"000012521";
		when x"00e75" => DOUT <= x"0000125a0";
		when x"00e76" => DOUT <= x"0002125c1";
		when x"00e77" => DOUT <= x"0002125c0";
		when x"00e78" => DOUT <= x"0000125a1";
		when x"00e79" => DOUT <= x"000012520";
		when x"00e7a" => DOUT <= x"000212541";
		when x"00e7b" => DOUT <= x"000212540";
		when x"00e7c" => DOUT <= x"000012521";
		when x"00e7d" => DOUT <= x"0000125a0";
		when x"00e7e" => DOUT <= x"0002125c1";
		when x"00e7f" => DOUT <= x"0002125c0";
		when x"00e80" => DOUT <= x"0000125a1";
		when x"00e81" => DOUT <= x"000012520";
		when x"00e82" => DOUT <= x"000212541";
		when x"00e83" => DOUT <= x"000212540";
		when x"00e84" => DOUT <= x"000012521";
		when x"00e85" => DOUT <= x"0000125a0";
		when x"00e86" => DOUT <= x"0002125c1";
		when x"00e87" => DOUT <= x"0002125c0";
		when x"00e88" => DOUT <= x"0000125a1";
		when x"00e89" => DOUT <= x"000012520";
		when x"00e8a" => DOUT <= x"000212541";
		when x"00e8b" => DOUT <= x"000212540";
		when x"00e8c" => DOUT <= x"000012521";
		when x"00e8d" => DOUT <= x"0000125a0";
		when x"00e8e" => DOUT <= x"0002125c1";
		when x"00e8f" => DOUT <= x"0002125c0";
		when x"00e90" => DOUT <= x"0000125a1";
		when x"00e91" => DOUT <= x"000012520";
		when x"00e92" => DOUT <= x"000212541";
		when x"00e93" => DOUT <= x"000212540";
		when x"00e94" => DOUT <= x"000012521";
		when x"00e95" => DOUT <= x"0000125a0";
		when x"00e96" => DOUT <= x"0002125c1";
		when x"00e97" => DOUT <= x"0002125c0";
		when x"00e98" => DOUT <= x"0000125a1";
		when x"00e99" => DOUT <= x"000012520";
		when x"00e9a" => DOUT <= x"000212541";
		when x"00e9b" => DOUT <= x"000212540";
		when x"00e9c" => DOUT <= x"000012521";
		when x"00e9d" => DOUT <= x"0000125a0";
		when x"00e9e" => DOUT <= x"0002125c1";
		when x"00e9f" => DOUT <= x"0002125c0";
		when x"00ea0" => DOUT <= x"0000125a1";
		when x"00ea1" => DOUT <= x"000012520";
		when x"00ea2" => DOUT <= x"000212541";
		when x"00ea3" => DOUT <= x"000212540";
		when x"00ea4" => DOUT <= x"000012521";
		when x"00ea5" => DOUT <= x"0000125a0";
		when x"00ea6" => DOUT <= x"0002125c1";
		when x"00ea7" => DOUT <= x"0002125c0";
		when x"00ea8" => DOUT <= x"0000125a1";
		when x"00ea9" => DOUT <= x"000012520";
		when x"00eaa" => DOUT <= x"000212541";
		when x"00eab" => DOUT <= x"000212540";
		when x"00eac" => DOUT <= x"000012521";
		when x"00ead" => DOUT <= x"0000125a0";
		when x"00eae" => DOUT <= x"0002125c1";
		when x"00eaf" => DOUT <= x"0002125c0";
		when x"00eb0" => DOUT <= x"0000021a1";
		when x"00eb1" => DOUT <= x"000002120";
		when x"00eb2" => DOUT <= x"000202141";
		when x"00eb3" => DOUT <= x"000202140";
		when x"00eb4" => DOUT <= x"000002121";
		when x"00eb5" => DOUT <= x"0000021a0";
		when x"00eb6" => DOUT <= x"0002021c1";
		when x"00eb7" => DOUT <= x"0002021c0";
		when x"00eb8" => DOUT <= x"0000021a1";
		when x"00eb9" => DOUT <= x"000002120";
		when x"00eba" => DOUT <= x"000202141";
		when x"00ebb" => DOUT <= x"000202140";
		when x"00ebc" => DOUT <= x"000002121";
		when x"00ebd" => DOUT <= x"0000021a0";
		when x"00ebe" => DOUT <= x"0002021c1";
		when x"00ebf" => DOUT <= x"0002021c0";
		when x"00ec0" => DOUT <= x"0000021a1";
		when x"00ec1" => DOUT <= x"000002120";
		when x"00ec2" => DOUT <= x"000202141";
		when x"00ec3" => DOUT <= x"000202140";
		when x"00ec4" => DOUT <= x"000002121";
		when x"00ec5" => DOUT <= x"0000021a0";
		when x"00ec6" => DOUT <= x"0002021c1";
		when x"00ec7" => DOUT <= x"0002021c0";
		when x"00ec8" => DOUT <= x"0000021a1";
		when x"00ec9" => DOUT <= x"000002120";
		when x"00eca" => DOUT <= x"000202141";
		when x"00ecb" => DOUT <= x"000202140";
		when x"00ecc" => DOUT <= x"000002121";
		when x"00ecd" => DOUT <= x"0000021a0";
		when x"00ece" => DOUT <= x"0002021c1";
		when x"00ecf" => DOUT <= x"0002021c0";
		when x"00ed0" => DOUT <= x"0000025a5";
		when x"00ed1" => DOUT <= x"000002524";
		when x"00ed2" => DOUT <= x"000202545";
		when x"00ed3" => DOUT <= x"000202544";
		when x"00ed4" => DOUT <= x"000002525";
		when x"00ed5" => DOUT <= x"0000025a4";
		when x"00ed6" => DOUT <= x"0002025c5";
		when x"00ed7" => DOUT <= x"0002025c4";
		when x"00ed8" => DOUT <= x"0000025a5";
		when x"00ed9" => DOUT <= x"000002524";
		when x"00eda" => DOUT <= x"000202545";
		when x"00edb" => DOUT <= x"000202544";
		when x"00edc" => DOUT <= x"000002525";
		when x"00edd" => DOUT <= x"0000025a4";
		when x"00ede" => DOUT <= x"0002025c5";
		when x"00edf" => DOUT <= x"0002025c4";
		when x"00ee0" => DOUT <= x"0000025a5";
		when x"00ee1" => DOUT <= x"000002524";
		when x"00ee2" => DOUT <= x"000202545";
		when x"00ee3" => DOUT <= x"000202544";
		when x"00ee4" => DOUT <= x"000002525";
		when x"00ee5" => DOUT <= x"0000025a4";
		when x"00ee6" => DOUT <= x"0002025c5";
		when x"00ee7" => DOUT <= x"0002025c4";
		when x"00ee8" => DOUT <= x"0000025a5";
		when x"00ee9" => DOUT <= x"000002524";
		when x"00eea" => DOUT <= x"000202545";
		when x"00eeb" => DOUT <= x"000202544";
		when x"00eec" => DOUT <= x"000002525";
		when x"00eed" => DOUT <= x"0000025a4";
		when x"00eee" => DOUT <= x"0002025c5";
		when x"00eef" => DOUT <= x"0002025c4";
		when x"00ef0" => DOUT <= x"0000027a5";
		when x"00ef1" => DOUT <= x"000002724";
		when x"00ef2" => DOUT <= x"000202745";
		when x"00ef3" => DOUT <= x"000202744";
		when x"00ef4" => DOUT <= x"000002725";
		when x"00ef5" => DOUT <= x"0000027a4";
		when x"00ef6" => DOUT <= x"0002027c5";
		when x"00ef7" => DOUT <= x"0002027c4";
		when x"00ef8" => DOUT <= x"0000127a5";
		when x"00ef9" => DOUT <= x"000012724";
		when x"00efa" => DOUT <= x"000212745";
		when x"00efb" => DOUT <= x"000202744";
		when x"00efc" => DOUT <= x"000002725";
		when x"00efd" => DOUT <= x"0000027a4";
		when x"00efe" => DOUT <= x"0002027c5";
		when x"00eff" => DOUT <= x"0002027c4";
		when x"00f00" => DOUT <= x"0000027a5";
		when x"00f01" => DOUT <= x"000002724";
		when x"00f02" => DOUT <= x"000202745";
		when x"00f03" => DOUT <= x"000202744";
		when x"00f04" => DOUT <= x"000002725";
		when x"00f05" => DOUT <= x"0000027a4";
		when x"00f06" => DOUT <= x"0002027c5";
		when x"00f07" => DOUT <= x"0002027c4";
		when x"00f08" => DOUT <= x"0000027a5";
		when x"00f09" => DOUT <= x"000002724";
		when x"00f0a" => DOUT <= x"000202745";
		when x"00f0b" => DOUT <= x"000202744";
		when x"00f0c" => DOUT <= x"000002725";
		when x"00f0d" => DOUT <= x"0000027a4";
		when x"00f0e" => DOUT <= x"0002027c5";
		when x"00f0f" => DOUT <= x"0002027c4";
		when x"00f10" => DOUT <= x"0000025a5";
		when x"00f11" => DOUT <= x"000002524";
		when x"00f12" => DOUT <= x"000202545";
		when x"00f13" => DOUT <= x"000202544";
		when x"00f14" => DOUT <= x"000002525";
		when x"00f15" => DOUT <= x"0000025a4";
		when x"00f16" => DOUT <= x"0002025c5";
		when x"00f17" => DOUT <= x"0002025c4";
		when x"00f18" => DOUT <= x"0000125a5";
		when x"00f19" => DOUT <= x"000012524";
		when x"00f1a" => DOUT <= x"000212545";
		when x"00f1b" => DOUT <= x"000202544";
		when x"00f1c" => DOUT <= x"000002525";
		when x"00f1d" => DOUT <= x"0000025a4";
		when x"00f1e" => DOUT <= x"0002025c5";
		when x"00f1f" => DOUT <= x"0002025c4";
		when x"00f20" => DOUT <= x"0000025a5";
		when x"00f21" => DOUT <= x"000002524";
		when x"00f22" => DOUT <= x"000202545";
		when x"00f23" => DOUT <= x"000202544";
		when x"00f24" => DOUT <= x"000002525";
		when x"00f25" => DOUT <= x"0000025a4";
		when x"00f26" => DOUT <= x"0002025c5";
		when x"00f27" => DOUT <= x"0002025c4";
		when x"00f28" => DOUT <= x"0000025a5";
		when x"00f29" => DOUT <= x"000002524";
		when x"00f2a" => DOUT <= x"000202545";
		when x"00f2b" => DOUT <= x"000202544";
		when x"00f2c" => DOUT <= x"000002525";
		when x"00f2d" => DOUT <= x"0000025a4";
		when x"00f2e" => DOUT <= x"0002025c5";
		when x"00f2f" => DOUT <= x"0002025c4";
		when x"00f30" => DOUT <= x"0000027a5";
		when x"00f31" => DOUT <= x"000002724";
		when x"00f32" => DOUT <= x"000202745";
		when x"00f33" => DOUT <= x"000202744";
		when x"00f34" => DOUT <= x"000002725";
		when x"00f35" => DOUT <= x"0000027a4";
		when x"00f36" => DOUT <= x"0002027c5";
		when x"00f37" => DOUT <= x"0002027c4";
		when x"00f38" => DOUT <= x"0000027a5";
		when x"00f39" => DOUT <= x"000002724";
		when x"00f3a" => DOUT <= x"000202745";
		when x"00f3b" => DOUT <= x"000202744";
		when x"00f3c" => DOUT <= x"000002725";
		when x"00f3d" => DOUT <= x"0000027a4";
		when x"00f3e" => DOUT <= x"0002027c5";
		when x"00f3f" => DOUT <= x"0002027c4";
		when x"00f40" => DOUT <= x"0000027a5";
		when x"00f41" => DOUT <= x"000002724";
		when x"00f42" => DOUT <= x"000202745";
		when x"00f43" => DOUT <= x"000202744";
		when x"00f44" => DOUT <= x"000002725";
		when x"00f45" => DOUT <= x"0000027a4";
		when x"00f46" => DOUT <= x"0002027c5";
		when x"00f47" => DOUT <= x"0002027c4";
		when x"00f48" => DOUT <= x"0000027a5";
		when x"00f49" => DOUT <= x"000002724";
		when x"00f4a" => DOUT <= x"000202745";
		when x"00f4b" => DOUT <= x"000202744";
		when x"00f4c" => DOUT <= x"000002725";
		when x"00f4d" => DOUT <= x"0000027a4";
		when x"00f4e" => DOUT <= x"0002027c5";
		when x"00f4f" => DOUT <= x"0002027c4";
		when x"00f50" => DOUT <= x"0000027a5";
		when x"00f51" => DOUT <= x"000002724";
		when x"00f52" => DOUT <= x"000202745";
		when x"00f53" => DOUT <= x"000202744";
		when x"00f54" => DOUT <= x"000002725";
		when x"00f55" => DOUT <= x"0000027a4";
		when x"00f56" => DOUT <= x"0002027c5";
		when x"00f57" => DOUT <= x"0002027c4";
		when x"00f58" => DOUT <= x"0000027a5";
		when x"00f59" => DOUT <= x"000002724";
		when x"00f5a" => DOUT <= x"000202745";
		when x"00f5b" => DOUT <= x"000202744";
		when x"00f5c" => DOUT <= x"000002725";
		when x"00f5d" => DOUT <= x"0000027a4";
		when x"00f5e" => DOUT <= x"0002027c5";
		when x"00f5f" => DOUT <= x"0002027c4";
		when x"00f60" => DOUT <= x"0000027a5";
		when x"00f61" => DOUT <= x"000002724";
		when x"00f62" => DOUT <= x"000202745";
		when x"00f63" => DOUT <= x"000202744";
		when x"00f64" => DOUT <= x"000002725";
		when x"00f65" => DOUT <= x"0000027a4";
		when x"00f66" => DOUT <= x"0002027c5";
		when x"00f67" => DOUT <= x"0002027c4";
		when x"00f68" => DOUT <= x"0000027a5";
		when x"00f69" => DOUT <= x"000002724";
		when x"00f6a" => DOUT <= x"000202745";
		when x"00f6b" => DOUT <= x"000202744";
		when x"00f6c" => DOUT <= x"000002725";
		when x"00f6d" => DOUT <= x"0000027a4";
		when x"00f6e" => DOUT <= x"0002027c5";
		when x"00f6f" => DOUT <= x"0002027c4";
		when x"00f70" => DOUT <= x"0000025a5";
		when x"00f71" => DOUT <= x"000002524";
		when x"00f72" => DOUT <= x"000202545";
		when x"00f73" => DOUT <= x"000202544";
		when x"00f74" => DOUT <= x"000002525";
		when x"00f75" => DOUT <= x"0000025a4";
		when x"00f76" => DOUT <= x"0002025c5";
		when x"00f77" => DOUT <= x"0002025c4";
		when x"00f78" => DOUT <= x"0000025a5";
		when x"00f79" => DOUT <= x"000002524";
		when x"00f7a" => DOUT <= x"000202545";
		when x"00f7b" => DOUT <= x"000202544";
		when x"00f7c" => DOUT <= x"000002525";
		when x"00f7d" => DOUT <= x"0000025a4";
		when x"00f7e" => DOUT <= x"0002025c5";
		when x"00f7f" => DOUT <= x"0002025c4";
		when x"00f80" => DOUT <= x"0000025a5";
		when x"00f81" => DOUT <= x"000002524";
		when x"00f82" => DOUT <= x"000202545";
		when x"00f83" => DOUT <= x"000202544";
		when x"00f84" => DOUT <= x"000002525";
		when x"00f85" => DOUT <= x"0000025a4";
		when x"00f86" => DOUT <= x"0002025c5";
		when x"00f87" => DOUT <= x"0002025c4";
		when x"00f88" => DOUT <= x"0000025a5";
		when x"00f89" => DOUT <= x"000002524";
		when x"00f8a" => DOUT <= x"000202545";
		when x"00f8b" => DOUT <= x"000202544";
		when x"00f8c" => DOUT <= x"000002525";
		when x"00f8d" => DOUT <= x"0000025a4";
		when x"00f8e" => DOUT <= x"0002025c5";
		when x"00f8f" => DOUT <= x"0002025c4";
		when x"00f90" => DOUT <= x"0000025a5";
		when x"00f91" => DOUT <= x"000002524";
		when x"00f92" => DOUT <= x"000202545";
		when x"00f93" => DOUT <= x"000202544";
		when x"00f94" => DOUT <= x"000002525";
		when x"00f95" => DOUT <= x"0000025a4";
		when x"00f96" => DOUT <= x"0002025c5";
		when x"00f97" => DOUT <= x"0002025c4";
		when x"00f98" => DOUT <= x"0000025a5";
		when x"00f99" => DOUT <= x"000002524";
		when x"00f9a" => DOUT <= x"000202545";
		when x"00f9b" => DOUT <= x"000202544";
		when x"00f9c" => DOUT <= x"000002525";
		when x"00f9d" => DOUT <= x"0000025a4";
		when x"00f9e" => DOUT <= x"0002025c5";
		when x"00f9f" => DOUT <= x"0002025c4";
		when x"00fa0" => DOUT <= x"0000025a5";
		when x"00fa1" => DOUT <= x"000002524";
		when x"00fa2" => DOUT <= x"000202545";
		when x"00fa3" => DOUT <= x"000202544";
		when x"00fa4" => DOUT <= x"000002525";
		when x"00fa5" => DOUT <= x"0000025a4";
		when x"00fa6" => DOUT <= x"0002025c5";
		when x"00fa7" => DOUT <= x"0002025c4";
		when x"00fa8" => DOUT <= x"0000025a5";
		when x"00fa9" => DOUT <= x"000002524";
		when x"00faa" => DOUT <= x"000202545";
		when x"00fab" => DOUT <= x"000202544";
		when x"00fac" => DOUT <= x"000002525";
		when x"00fad" => DOUT <= x"0000025a4";
		when x"00fae" => DOUT <= x"0002025c5";
		when x"00faf" => DOUT <= x"0002025c4";
		when x"00fb0" => DOUT <= x"0000021a1";
		when x"00fb1" => DOUT <= x"000002120";
		when x"00fb2" => DOUT <= x"000202141";
		when x"00fb3" => DOUT <= x"000202140";
		when x"00fb4" => DOUT <= x"000002121";
		when x"00fb5" => DOUT <= x"0000021a0";
		when x"00fb6" => DOUT <= x"0002021c1";
		when x"00fb7" => DOUT <= x"0002021c0";
		when x"00fb8" => DOUT <= x"0000021a1";
		when x"00fb9" => DOUT <= x"000002120";
		when x"00fba" => DOUT <= x"000202141";
		when x"00fbb" => DOUT <= x"000202140";
		when x"00fbc" => DOUT <= x"000002121";
		when x"00fbd" => DOUT <= x"0000021a0";
		when x"00fbe" => DOUT <= x"0002021c1";
		when x"00fbf" => DOUT <= x"0002021c0";
		when x"00fc0" => DOUT <= x"0000021a1";
		when x"00fc1" => DOUT <= x"000002120";
		when x"00fc2" => DOUT <= x"000202141";
		when x"00fc3" => DOUT <= x"000202140";
		when x"00fc4" => DOUT <= x"000002121";
		when x"00fc5" => DOUT <= x"0000021a0";
		when x"00fc6" => DOUT <= x"0002021c1";
		when x"00fc7" => DOUT <= x"0002021c0";
		when x"00fc8" => DOUT <= x"0000021a1";
		when x"00fc9" => DOUT <= x"000002120";
		when x"00fca" => DOUT <= x"000202141";
		when x"00fcb" => DOUT <= x"000202140";
		when x"00fcc" => DOUT <= x"000002121";
		when x"00fcd" => DOUT <= x"0000021a0";
		when x"00fce" => DOUT <= x"0002021c1";
		when x"00fcf" => DOUT <= x"0002021c0";
		when x"00fd0" => DOUT <= x"000002901";
		when x"00fd1" => DOUT <= x"000002900";
		when x"00fd2" => DOUT <= x"000002901";
		when x"00fd3" => DOUT <= x"000002900";
		when x"00fd4" => DOUT <= x"000002181";
		when x"00fd5" => DOUT <= x"000002100";
		when x"00fd6" => DOUT <= x"000002101";
		when x"00fd7" => DOUT <= x"000002100";
		when x"00fd8" => DOUT <= x"000002101";
		when x"00fd9" => DOUT <= x"000002180";
		when x"00fda" => DOUT <= x"000002181";
		when x"00fdb" => DOUT <= x"000002180";
		when x"00fdc" => DOUT <= x"000002181";
		when x"00fdd" => DOUT <= x"000002100";
		when x"00fde" => DOUT <= x"000002101";
		when x"00fdf" => DOUT <= x"000002100";
		when x"00fe0" => DOUT <= x"000002101";
		when x"00fe1" => DOUT <= x"000002180";
		when x"00fe2" => DOUT <= x"000002181";
		when x"00fe3" => DOUT <= x"000002180";
          when others => 
    end case;
end if;

end process;

end behavior;
