library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

---- Uncomment the following library declaration if instantiating
---- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity instrom is
    Port ( CLK : in std_logic;
           ADDR : in std_logic_vector(18 DOWNTO 0);
           DOUT : out std_logic_vector(35 DOWNTO 0)
           );
end instrom;


architecture behavior of instrom is

begin

main: Process(CLK)
begin
If (falling_edge(CLK)) Then
    case ADDR is

		when b"0000000000000000000" => DOUT <= x"010000fd0";
		when b"0000000000000000001" => DOUT <= x"028fffff6";
		when b"0000000000000000010" => DOUT <= x"010000fd0";
		when b"0000000000000000011" => DOUT <= x"00c000000";
		when b"0000000000000000100" => DOUT <= x"088000002";
		when b"0000000000000000101" => DOUT <= x"010000fd4";
		when b"0000000000000000110" => DOUT <= x"028fffff5";
		when b"0000000000000000111" => DOUT <= x"0e8fffffd";
		when b"0000000000000001000" => DOUT <= x"208000000";
		when b"0000000000000001001" => DOUT <= x"108000008";
		when b"0000000000000001010" => DOUT <= x"07800000f";
		when b"0000000000000001011" => DOUT <= x"010000fd4";
		when b"0000000000000001100" => DOUT <= x"0e8fffffc";
		when b"0000000000000001101" => DOUT <= x"208000000";
		when b"0000000000000001110" => DOUT <= x"10800000d";
		when b"0000000000000001111" => DOUT <= x"010000fd4";
		when b"0000000000000010000" => DOUT <= x"038fffffe";
		when b"0000000000000010001" => DOUT <= x"0e8fffffd";
		when b"0000000000000010010" => DOUT <= x"008000000";
		when b"0000000000000010011" => DOUT <= x"208000000";
		when b"0000000000000010100" => DOUT <= x"108000013";
		when b"0000000000000010101" => DOUT <= x"010000fd4";
		when b"0000000000000010110" => DOUT <= x"0e8fffffd";
		when b"0000000000000010111" => DOUT <= x"208000000";
		when b"0000000000000011000" => DOUT <= x"108000017";
		when b"0000000000000011001" => DOUT <= x"00a000000";
		when b"0000000000000011010" => DOUT <= x"098000015";
		when b"0000000000000011011" => DOUT <= x"010000fd4";
		when b"0000000000000011100" => DOUT <= x"0e8fffffd";
		when b"0000000000000011101" => DOUT <= x"208000000";
		when b"0000000000000011110" => DOUT <= x"10800001d";
		when b"0000000000000011111" => DOUT <= x"00c000000";
		when b"0000000000000100000" => DOUT <= x"08800000b";
		when b"0000000000000100001" => DOUT <= x"010000fb0";
		when b"0000000000000100010" => DOUT <= x"028fffffc";
		when b"0000000000000100011" => DOUT <= x"0e8fffff9";
		when b"0000000000000100100" => DOUT <= x"008000000";
		when b"0000000000000100101" => DOUT <= x"208000000";
		when b"0000000000000100110" => DOUT <= x"108000025";
		when b"0000000000000100111" => DOUT <= x"010000fb0";
		when b"0000000000000101000" => DOUT <= x"0e8fffff9";
		when b"0000000000000101001" => DOUT <= x"208000000";
		when b"0000000000000101010" => DOUT <= x"108000029";
		when b"0000000000000101011" => DOUT <= x"00c000000";
		when b"0000000000000101100" => DOUT <= x"088000027";
		when b"0000000000000101101" => DOUT <= x"010000000";
		when b"0000000000000101110" => DOUT <= x"0e8fffffc";
		when b"0000000000000101111" => DOUT <= x"208000000";
		when b"0000000000000110000" => DOUT <= x"10800002f";
		when b"0000000000000110001" => DOUT <= x"010000010";
		when b"0000000000000110010" => DOUT <= x"0e8ffff18";
		when b"0000000000000110011" => DOUT <= x"208000000";
		when b"0000000000000110100" => DOUT <= x"108000033";
		when b"0000000000000110101" => DOUT <= x"0100003b0";
		when b"0000000000000110110" => DOUT <= x"0e8ffff30";
		when b"0000000000000110111" => DOUT <= x"208000000";
		when b"0000000000000111000" => DOUT <= x"108000037";
		when b"0000000000000111001" => DOUT <= x"0100006f0";
		when b"0000000000000111010" => DOUT <= x"0e8ffff30";
		when b"0000000000000111011" => DOUT <= x"208000000";
		when b"0000000000000111100" => DOUT <= x"10800003b";
		when b"0000000000000111101" => DOUT <= x"010000a30";
		when b"0000000000000111110" => DOUT <= x"0e8ffff30";
		when b"0000000000000111111" => DOUT <= x"208000000";
		when b"0000000000001000000" => DOUT <= x"10800003f";
		when b"0000000000001000001" => DOUT <= x"010000000";
		when b"0000000000001000010" => DOUT <= x"0e8fffffc";
		when b"0000000000001000011" => DOUT <= x"208000000";
		when b"0000000000001000100" => DOUT <= x"108000043";
		when b"0000000000001000101" => DOUT <= x"010000dc0";
		when b"0000000000001000110" => DOUT <= x"028fffff4";
		when b"0000000000001000111" => DOUT <= x"0e8fffff9";
		when b"0000000000001001000" => DOUT <= x"008000000";
		when b"0000000000001001001" => DOUT <= x"208000000";
		when b"0000000000001001010" => DOUT <= x"108000049";
		when b"0000000000001001011" => DOUT <= x"010000dc0";
		when b"0000000000001001100" => DOUT <= x"0e8fffff9";
		when b"0000000000001001101" => DOUT <= x"208000000";
		when b"0000000000001001110" => DOUT <= x"10800004d";
		when b"0000000000001001111" => DOUT <= x"00c000000";
		when b"0000000000001010000" => DOUT <= x"08800004b";
		when b"0000000000001010001" => DOUT <= x"010000de0";
		when b"0000000000001010010" => DOUT <= x"0e8fffff8";
		when b"0000000000001010011" => DOUT <= x"208000000";
		when b"0000000000001010100" => DOUT <= x"108000053";
		when b"0000000000001010101" => DOUT <= x"010000e00";
		when b"0000000000001010110" => DOUT <= x"028ffff50";
		when b"0000000000001010111" => DOUT <= x"0e8fffff9";
		when b"0000000000001011000" => DOUT <= x"008000000";
		when b"0000000000001011001" => DOUT <= x"208000000";
		when b"0000000000001011010" => DOUT <= x"108000059";
		when b"0000000000001011011" => DOUT <= x"010000e00";
		when b"0000000000001011100" => DOUT <= x"0e8fffff9";
		when b"0000000000001011101" => DOUT <= x"208000000";
		when b"0000000000001011110" => DOUT <= x"10800005d";
		when b"0000000000001011111" => DOUT <= x"00c000000";
		when b"0000000000001100000" => DOUT <= x"08800005b";
		when b"0000000000001100001" => DOUT <= x"010000e30";
		when b"0000000000001100010" => DOUT <= x"028ffff38";
		when b"0000000000001100011" => DOUT <= x"0e8fffff9";
		when b"0000000000001100100" => DOUT <= x"008000000";
		when b"0000000000001100101" => DOUT <= x"208000000";
		when b"0000000000001100110" => DOUT <= x"108000065";
		when b"0000000000001100111" => DOUT <= x"010000e30";
		when b"0000000000001101000" => DOUT <= x"0e8fffff9";
		when b"0000000000001101001" => DOUT <= x"208000000";
		when b"0000000000001101010" => DOUT <= x"108000069";
		when b"0000000000001101011" => DOUT <= x"00c000000";
		when b"0000000000001101100" => DOUT <= x"088000067";
		when b"0000000000001101101" => DOUT <= x"010000e50";
		when b"0000000000001101110" => DOUT <= x"028fffd80";
		when b"0000000000001101111" => DOUT <= x"0e8fffff9";
		when b"0000000000001110000" => DOUT <= x"008000000";
		when b"0000000000001110001" => DOUT <= x"208000000";
		when b"0000000000001110010" => DOUT <= x"108000071";
		when b"0000000000001110011" => DOUT <= x"010000e50";
		when b"0000000000001110100" => DOUT <= x"0e8fffff9";
		when b"0000000000001110101" => DOUT <= x"208000000";
		when b"0000000000001110110" => DOUT <= x"108000075";
		when b"0000000000001110111" => DOUT <= x"00c000000";
		when b"0000000000001111000" => DOUT <= x"088000073";
		when b"0000000000001111001" => DOUT <= x"010000e70";
		when b"0000000000001111010" => DOUT <= x"028ffffec";
		when b"0000000000001111011" => DOUT <= x"0e8fffff9";
		when b"0000000000001111100" => DOUT <= x"008000000";
		when b"0000000000001111101" => DOUT <= x"208000000";
		when b"0000000000001111110" => DOUT <= x"10800007d";
		when b"0000000000001111111" => DOUT <= x"010000e70";
		when b"0000000000010000000" => DOUT <= x"0e8fffff9";
		when b"0000000000010000001" => DOUT <= x"208000000";
		when b"0000000000010000010" => DOUT <= x"108000081";
		when b"0000000000010000011" => DOUT <= x"00c000000";
		when b"0000000000010000100" => DOUT <= x"08800007f";
		when b"0000000000010000101" => DOUT <= x"010000f30";
		when b"0000000000010000110" => DOUT <= x"028fffdf7";
		when b"0000000000010000111" => DOUT <= x"0e8fffff9";
		when b"0000000000010001000" => DOUT <= x"208000000";
		when b"0000000000010001001" => DOUT <= x"108000088";
		when b"0000000000010001010" => DOUT <= x"07800008f";
		when b"0000000000010001011" => DOUT <= x"010000f30";
		when b"0000000000010001100" => DOUT <= x"0e8fffff8";
		when b"0000000000010001101" => DOUT <= x"208000000";
		when b"0000000000010001110" => DOUT <= x"10800008d";
		when b"0000000000010001111" => DOUT <= x"010000f30";
		when b"0000000000010010000" => DOUT <= x"0e8fffff8";
		when b"0000000000010010001" => DOUT <= x"208000000";
		when b"0000000000010010010" => DOUT <= x"108000091";
		when b"0000000000010010011" => DOUT <= x"010000f50";
		when b"0000000000010010100" => DOUT <= x"038ffffec";
		when b"0000000000010010101" => DOUT <= x"0e8fffff9";
		when b"0000000000010010110" => DOUT <= x"008000000";
		when b"0000000000010010111" => DOUT <= x"208000000";
		when b"0000000000010011000" => DOUT <= x"108000097";
		when b"0000000000010011001" => DOUT <= x"010000f50";
		when b"0000000000010011010" => DOUT <= x"0e8fffff9";
		when b"0000000000010011011" => DOUT <= x"208000000";
		when b"0000000000010011100" => DOUT <= x"10800009b";
		when b"0000000000010011101" => DOUT <= x"00a000000";
		when b"0000000000010011110" => DOUT <= x"098000099";
		when b"0000000000010011111" => DOUT <= x"010000f70";
		when b"0000000000010100000" => DOUT <= x"038fffff6";
		when b"0000000000010100001" => DOUT <= x"0e8fffff9";
		when b"0000000000010100010" => DOUT <= x"008000000";
		when b"0000000000010100011" => DOUT <= x"208000000";
		when b"0000000000010100100" => DOUT <= x"1080000a3";
		when b"0000000000010100101" => DOUT <= x"010000f70";
		when b"0000000000010100110" => DOUT <= x"0e8fffff9";
		when b"0000000000010100111" => DOUT <= x"208000000";
		when b"0000000000010101000" => DOUT <= x"1080000a7";
		when b"0000000000010101001" => DOUT <= x"00a000000";
		when b"0000000000010101010" => DOUT <= x"0980000a5";
		when b"0000000000010101011" => DOUT <= x"010000f10";
		when b"0000000000010101100" => DOUT <= x"0e8fffff8";
		when b"0000000000010101101" => DOUT <= x"208000000";
		when b"0000000000010101110" => DOUT <= x"1080000ad";
		when b"0000000000010101111" => DOUT <= x"010000f70";
		when b"0000000000010110000" => DOUT <= x"038fffff7";
		when b"0000000000010110001" => DOUT <= x"0e8fffff9";
		when b"0000000000010110010" => DOUT <= x"008000000";
		when b"0000000000010110011" => DOUT <= x"208000000";
		when b"0000000000010110100" => DOUT <= x"1080000b3";
		when b"0000000000010110101" => DOUT <= x"010000f70";
		when b"0000000000010110110" => DOUT <= x"0e8fffff9";
		when b"0000000000010110111" => DOUT <= x"208000000";
		when b"0000000000010111000" => DOUT <= x"1080000b7";
		when b"0000000000010111001" => DOUT <= x"00a000000";
		when b"0000000000010111010" => DOUT <= x"0980000b5";
		when b"0000000000010111011" => DOUT <= x"010000f90";
		when b"0000000000010111100" => DOUT <= x"0e8fffff9";
		when b"0000000000010111101" => DOUT <= x"208000000";
		when b"0000000000010111110" => DOUT <= x"1080000bd";
		when b"0000000000010111111" => DOUT <= x"00c000000";
		when b"0000000000011000000" => DOUT <= x"08800008b";
		when b"0000000000011000001" => DOUT <= x"010000fb0";
		when b"0000000000011000010" => DOUT <= x"028fffffc";
		when b"0000000000011000011" => DOUT <= x"0e8fffff9";
		when b"0000000000011000100" => DOUT <= x"008000000";
		when b"0000000000011000101" => DOUT <= x"208000000";
		when b"0000000000011000110" => DOUT <= x"1080000c5";
		when b"0000000000011000111" => DOUT <= x"010000fb0";
		when b"0000000000011001000" => DOUT <= x"0e8fffff9";
		when b"0000000000011001001" => DOUT <= x"208000000";
		when b"0000000000011001010" => DOUT <= x"1080000c9";
		when b"0000000000011001011" => DOUT <= x"00c000000";
		when b"0000000000011001100" => DOUT <= x"0880000c7";
		when b"0000000000011001101" => DOUT <= x"010000d70";
		when b"0000000000011001110" => DOUT <= x"0e8fffffc";
		when b"0000000000011001111" => DOUT <= x"208000000";
		when b"0000000000011010000" => DOUT <= x"1080000cf";
		when b"0000000000011010001" => DOUT <= x"010000d80";
		when b"0000000000011010010" => DOUT <= x"028fffffe";
		when b"0000000000011010011" => DOUT <= x"0e8fffffd";
		when b"0000000000011010100" => DOUT <= x"008000000";
		when b"0000000000011010101" => DOUT <= x"208000000";
		when b"0000000000011010110" => DOUT <= x"1080000d5";
		when b"0000000000011010111" => DOUT <= x"010000d80";
		when b"0000000000011011000" => DOUT <= x"0e8fffffd";
		when b"0000000000011011001" => DOUT <= x"208000000";
		when b"0000000000011011010" => DOUT <= x"1080000d9";
		when b"0000000000011011011" => DOUT <= x"00c000000";
		when b"0000000000011011100" => DOUT <= x"0880000d7";
		when b"0000000000011011101" => DOUT <= x"010000d90";
		when b"0000000000011011110" => DOUT <= x"028fffefe";
		when b"0000000000011011111" => DOUT <= x"0e8fffffd";
		when b"0000000000011100000" => DOUT <= x"008000000";
		when b"0000000000011100001" => DOUT <= x"208000000";
		when b"0000000000011100010" => DOUT <= x"1080000e1";
		when b"0000000000011100011" => DOUT <= x"010000d90";
		when b"0000000000011100100" => DOUT <= x"0e8fffffd";
		when b"0000000000011100101" => DOUT <= x"208000000";
		when b"0000000000011100110" => DOUT <= x"1080000e5";
		when b"0000000000011100111" => DOUT <= x"00c000000";
		when b"0000000000011101000" => DOUT <= x"0880000e3";
		when b"0000000000011101001" => DOUT <= x"010000da0";
		when b"0000000000011101010" => DOUT <= x"028fffefc";
		when b"0000000000011101011" => DOUT <= x"0e8fffffd";
		when b"0000000000011101100" => DOUT <= x"008000000";
		when b"0000000000011101101" => DOUT <= x"208000000";
		when b"0000000000011101110" => DOUT <= x"1080000ed";
		when b"0000000000011101111" => DOUT <= x"010000da0";
		when b"0000000000011110000" => DOUT <= x"0e8fffffd";
		when b"0000000000011110001" => DOUT <= x"208000000";
		when b"0000000000011110010" => DOUT <= x"1080000f1";
		when b"0000000000011110011" => DOUT <= x"00c000000";
		when b"0000000000011110100" => DOUT <= x"0880000ef";
		when b"0000000000011110101" => DOUT <= x"010000db0";
		when b"0000000000011110110" => DOUT <= x"0e8fffffc";
		when b"0000000000011110111" => DOUT <= x"208000000";
		when b"0000000000011111000" => DOUT <= x"1080000f7";
		when b"0000000000011111001" => DOUT <= x"010000dc0";
		when b"0000000000011111010" => DOUT <= x"028fffff4";
		when b"0000000000011111011" => DOUT <= x"0e8fffff9";
		when b"0000000000011111100" => DOUT <= x"008000000";
		when b"0000000000011111101" => DOUT <= x"208000000";
		when b"0000000000011111110" => DOUT <= x"1080000fd";
		when b"0000000000011111111" => DOUT <= x"010000dc0";
		when b"0000000000100000000" => DOUT <= x"0e8fffff9";
		when b"0000000000100000001" => DOUT <= x"208000000";
		when b"0000000000100000010" => DOUT <= x"108000101";
		when b"0000000000100000011" => DOUT <= x"00c000000";
		when b"0000000000100000100" => DOUT <= x"0880000ff";
		when b"0000000000100000101" => DOUT <= x"010000de0";
		when b"0000000000100000110" => DOUT <= x"0e8fffff8";
		when b"0000000000100000111" => DOUT <= x"208000000";
		when b"0000000000100001000" => DOUT <= x"108000107";
		when b"0000000000100001001" => DOUT <= x"010000e00";
		when b"0000000000100001010" => DOUT <= x"028ffffe9";
		when b"0000000000100001011" => DOUT <= x"0e8fffff9";
		when b"0000000000100001100" => DOUT <= x"008000000";
		when b"0000000000100001101" => DOUT <= x"208000000";
		when b"0000000000100001110" => DOUT <= x"10800010d";
		when b"0000000000100001111" => DOUT <= x"010000e00";
		when b"0000000000100010000" => DOUT <= x"0e8fffff9";
		when b"0000000000100010001" => DOUT <= x"208000000";
		when b"0000000000100010010" => DOUT <= x"108000111";
		when b"0000000000100010011" => DOUT <= x"00c000000";
		when b"0000000000100010100" => DOUT <= x"08800010f";
		when b"0000000000100010101" => DOUT <= x"010000e30";
		when b"0000000000100010110" => DOUT <= x"028ffff38";
		when b"0000000000100010111" => DOUT <= x"0e8fffff9";
		when b"0000000000100011000" => DOUT <= x"008000000";
		when b"0000000000100011001" => DOUT <= x"208000000";
		when b"0000000000100011010" => DOUT <= x"108000119";
		when b"0000000000100011011" => DOUT <= x"010000e30";
		when b"0000000000100011100" => DOUT <= x"0e8fffff9";
		when b"0000000000100011101" => DOUT <= x"208000000";
		when b"0000000000100011110" => DOUT <= x"10800011d";
		when b"0000000000100011111" => DOUT <= x"00c000000";
		when b"0000000000100100000" => DOUT <= x"08800011b";
		when b"0000000000100100001" => DOUT <= x"010000e50";
		when b"0000000000100100010" => DOUT <= x"028fffd80";
		when b"0000000000100100011" => DOUT <= x"0e8fffff9";
		when b"0000000000100100100" => DOUT <= x"008000000";
		when b"0000000000100100101" => DOUT <= x"208000000";
		when b"0000000000100100110" => DOUT <= x"108000125";
		when b"0000000000100100111" => DOUT <= x"010000e50";
		when b"0000000000100101000" => DOUT <= x"0e8fffff9";
		when b"0000000000100101001" => DOUT <= x"208000000";
		when b"0000000000100101010" => DOUT <= x"108000129";
		when b"0000000000100101011" => DOUT <= x"00c000000";
		when b"0000000000100101100" => DOUT <= x"088000127";
		when b"0000000000100101101" => DOUT <= x"010000e70";
		when b"0000000000100101110" => DOUT <= x"028ffffec";
		when b"0000000000100101111" => DOUT <= x"0e8fffff9";
		when b"0000000000100110000" => DOUT <= x"008000000";
		when b"0000000000100110001" => DOUT <= x"208000000";
		when b"0000000000100110010" => DOUT <= x"108000131";
		when b"0000000000100110011" => DOUT <= x"010000e70";
		when b"0000000000100110100" => DOUT <= x"0e8fffff9";
		when b"0000000000100110101" => DOUT <= x"208000000";
		when b"0000000000100110110" => DOUT <= x"108000135";
		when b"0000000000100110111" => DOUT <= x"00c000000";
		when b"0000000000100111000" => DOUT <= x"088000133";
		when b"0000000000100111001" => DOUT <= x"010000f30";
		when b"0000000000100111010" => DOUT <= x"028fffdf8";
		when b"0000000000100111011" => DOUT <= x"0e8fffff9";
		when b"0000000000100111100" => DOUT <= x"208000000";
		when b"0000000000100111101" => DOUT <= x"10800013c";
		when b"0000000000100111110" => DOUT <= x"078000143";
		when b"0000000000100111111" => DOUT <= x"010000f30";
		when b"0000000000101000000" => DOUT <= x"0e8fffff8";
		when b"0000000000101000001" => DOUT <= x"208000000";
		when b"0000000000101000010" => DOUT <= x"108000141";
		when b"0000000000101000011" => DOUT <= x"010000f30";
		when b"0000000000101000100" => DOUT <= x"0e8fffff8";
		when b"0000000000101000101" => DOUT <= x"208000000";
		when b"0000000000101000110" => DOUT <= x"108000145";
		when b"0000000000101000111" => DOUT <= x"010000f50";
		when b"0000000000101001000" => DOUT <= x"038ffffec";
		when b"0000000000101001001" => DOUT <= x"0e8fffff9";
		when b"0000000000101001010" => DOUT <= x"008000000";
		when b"0000000000101001011" => DOUT <= x"208000000";
		when b"0000000000101001100" => DOUT <= x"10800014b";
		when b"0000000000101001101" => DOUT <= x"010000f50";
		when b"0000000000101001110" => DOUT <= x"0e8fffff9";
		when b"0000000000101001111" => DOUT <= x"208000000";
		when b"0000000000101010000" => DOUT <= x"10800014f";
		when b"0000000000101010001" => DOUT <= x"00a000000";
		when b"0000000000101010010" => DOUT <= x"09800014d";
		when b"0000000000101010011" => DOUT <= x"010000f70";
		when b"0000000000101010100" => DOUT <= x"038fffff6";
		when b"0000000000101010101" => DOUT <= x"0e8fffff9";
		when b"0000000000101010110" => DOUT <= x"008000000";
		when b"0000000000101010111" => DOUT <= x"208000000";
		when b"0000000000101011000" => DOUT <= x"108000157";
		when b"0000000000101011001" => DOUT <= x"010000f70";
		when b"0000000000101011010" => DOUT <= x"0e8fffff9";
		when b"0000000000101011011" => DOUT <= x"208000000";
		when b"0000000000101011100" => DOUT <= x"10800015b";
		when b"0000000000101011101" => DOUT <= x"00a000000";
		when b"0000000000101011110" => DOUT <= x"098000159";
		when b"0000000000101011111" => DOUT <= x"010000f10";
		when b"0000000000101100000" => DOUT <= x"0e8fffff8";
		when b"0000000000101100001" => DOUT <= x"208000000";
		when b"0000000000101100010" => DOUT <= x"108000161";
		when b"0000000000101100011" => DOUT <= x"010000f70";
		when b"0000000000101100100" => DOUT <= x"038fffff7";
		when b"0000000000101100101" => DOUT <= x"0e8fffff9";
		when b"0000000000101100110" => DOUT <= x"008000000";
		when b"0000000000101100111" => DOUT <= x"208000000";
		when b"0000000000101101000" => DOUT <= x"108000167";
		when b"0000000000101101001" => DOUT <= x"010000f70";
		when b"0000000000101101010" => DOUT <= x"0e8fffff9";
		when b"0000000000101101011" => DOUT <= x"208000000";
		when b"0000000000101101100" => DOUT <= x"10800016b";
		when b"0000000000101101101" => DOUT <= x"00a000000";
		when b"0000000000101101110" => DOUT <= x"098000169";
		when b"0000000000101101111" => DOUT <= x"010000f90";
		when b"0000000000101110000" => DOUT <= x"0e8fffff9";
		when b"0000000000101110001" => DOUT <= x"208000000";
		when b"0000000000101110010" => DOUT <= x"108000171";
		when b"0000000000101110011" => DOUT <= x"00c000000";
		when b"0000000000101110100" => DOUT <= x"08800013f";
		when b"0000000000101110101" => DOUT <= x"010000f30";
		when b"0000000000101110110" => DOUT <= x"0e8fffff8";
		when b"0000000000101110111" => DOUT <= x"208000000";
		when b"0000000000101111000" => DOUT <= x"108000177";
		when b"0000000000101111001" => DOUT <= x"010000f30";
		when b"0000000000101111010" => DOUT <= x"0e8fffff8";
		when b"0000000000101111011" => DOUT <= x"208000000";
		when b"0000000000101111100" => DOUT <= x"10800017b";
		when b"0000000000101111101" => DOUT <= x"010000f50";
		when b"0000000000101111110" => DOUT <= x"028ffffec";
		when b"0000000000101111111" => DOUT <= x"0e8fffff9";
		when b"0000000000110000000" => DOUT <= x"008000000";
		when b"0000000000110000001" => DOUT <= x"208000000";
		when b"0000000000110000010" => DOUT <= x"108000181";
		when b"0000000000110000011" => DOUT <= x"010000f50";
		when b"0000000000110000100" => DOUT <= x"0e8fffff9";
		when b"0000000000110000101" => DOUT <= x"208000000";
		when b"0000000000110000110" => DOUT <= x"108000185";
		when b"0000000000110000111" => DOUT <= x"00c000000";
		when b"0000000000110001000" => DOUT <= x"088000183";
		when b"0000000000110001001" => DOUT <= x"010000f70";
		when b"0000000000110001010" => DOUT <= x"028fffff6";
		when b"0000000000110001011" => DOUT <= x"0e8fffff9";
		when b"0000000000110001100" => DOUT <= x"008000000";
		when b"0000000000110001101" => DOUT <= x"208000000";
		when b"0000000000110001110" => DOUT <= x"10800018d";
		when b"0000000000110001111" => DOUT <= x"010000f70";
		when b"0000000000110010000" => DOUT <= x"0e8fffff9";
		when b"0000000000110010001" => DOUT <= x"208000000";
		when b"0000000000110010010" => DOUT <= x"108000191";
		when b"0000000000110010011" => DOUT <= x"00c000000";
		when b"0000000000110010100" => DOUT <= x"08800018f";
		when b"0000000000110010101" => DOUT <= x"010000f10";
		when b"0000000000110010110" => DOUT <= x"0e8fffff8";
		when b"0000000000110010111" => DOUT <= x"208000000";
		when b"0000000000110011000" => DOUT <= x"108000197";
		when b"0000000000110011001" => DOUT <= x"010000f70";
		when b"0000000000110011010" => DOUT <= x"028fffff7";
		when b"0000000000110011011" => DOUT <= x"0e8fffff9";
		when b"0000000000110011100" => DOUT <= x"008000000";
		when b"0000000000110011101" => DOUT <= x"208000000";
		when b"0000000000110011110" => DOUT <= x"10800019d";
		when b"0000000000110011111" => DOUT <= x"010000f70";
		when b"0000000000110100000" => DOUT <= x"0e8fffff9";
		when b"0000000000110100001" => DOUT <= x"208000000";
		when b"0000000000110100010" => DOUT <= x"1080001a1";
		when b"0000000000110100011" => DOUT <= x"00c000000";
		when b"0000000000110100100" => DOUT <= x"08800019f";
		when b"0000000000110100101" => DOUT <= x"010000f90";
		when b"0000000000110100110" => DOUT <= x"0e8fffff9";
		when b"0000000000110100111" => DOUT <= x"008000000";
		when b"0000000000110101000" => DOUT <= x"208000000";
		when b"0000000000110101001" => DOUT <= x"1080001a8";
		when b"0000000000110101010" => DOUT <= x"078000021";
			 when others =>
    end case;
end if;

end process;

end behavior;
